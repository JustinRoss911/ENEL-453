 fsd