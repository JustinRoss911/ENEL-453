library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_buzzing_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant d2buzz_LUT : array_1d := (

(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	0	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	995	)	,
(	1000	)	,
(	1005	)	,
(	1009	)	,
(	1014	)	,
(	1018	)	,
(	1023	)	,
(	1028	)	,
(	1032	)	,
(	1037	)	,
(	1041	)	,
(	1046	)	,
(	1051	)	,
(	1055	)	,
(	1060	)	,
(	1064	)	,
(	1069	)	,
(	1073	)	,
(	1078	)	,
(	1082	)	,
(	1087	)	,
(	1091	)	,
(	1096	)	,
(	1100	)	,
(	1105	)	,
(	1109	)	,
(	1113	)	,
(	1118	)	,
(	1122	)	,
(	1127	)	,
(	1131	)	,
(	1135	)	,
(	1140	)	,
(	1144	)	,
(	1148	)	,
(	1153	)	,
(	1157	)	,
(	1161	)	,
(	1166	)	,
(	1170	)	,
(	1174	)	,
(	1179	)	,
(	1183	)	,
(	1187	)	,
(	1191	)	,
(	1196	)	,
(	1200	)	,
(	1204	)	,
(	1208	)	,
(	1213	)	,
(	1217	)	,
(	1221	)	,
(	1225	)	,
(	1229	)	,
(	1234	)	,
(	1238	)	,
(	1242	)	,
(	1246	)	,
(	1250	)	,
(	1254	)	,
(	1259	)	,
(	1263	)	,
(	1267	)	,
(	1271	)	,
(	1275	)	,
(	1279	)	,
(	1283	)	,
(	1287	)	,
(	1291	)	,
(	1295	)	,
(	1299	)	,
(	1303	)	,
(	1307	)	,
(	1311	)	,
(	1315	)	,
(	1320	)	,
(	1324	)	,
(	1328	)	,
(	1332	)	,
(	1335	)	,
(	1339	)	,
(	1343	)	,
(	1347	)	,
(	1351	)	,
(	1355	)	,
(	1359	)	,
(	1363	)	,
(	1367	)	,
(	1371	)	,
(	1375	)	,
(	1379	)	,
(	1383	)	,
(	1387	)	,
(	1390	)	,
(	1394	)	,
(	1398	)	,
(	1402	)	,
(	1406	)	,
(	1410	)	,
(	1414	)	,
(	1417	)	,
(	1421	)	,
(	1425	)	,
(	1429	)	,
(	1433	)	,
(	1436	)	,
(	1440	)	,
(	1444	)	,
(	1448	)	,
(	1452	)	,
(	1455	)	,
(	1459	)	,
(	1463	)	,
(	1467	)	,
(	1470	)	,
(	1474	)	,
(	1478	)	,
(	1482	)	,
(	1485	)	,
(	1489	)	,
(	1493	)	,
(	1496	)	,
(	1500	)	,
(	1504	)	,
(	1507	)	,
(	1511	)	,
(	1515	)	,
(	1518	)	,
(	1522	)	,
(	1526	)	,
(	1529	)	,
(	1533	)	,
(	1537	)	,
(	1540	)	,
(	1544	)	,
(	1547	)	,
(	1551	)	,
(	1555	)	,
(	1558	)	,
(	1562	)	,
(	1565	)	,
(	1569	)	,
(	1572	)	,
(	1576	)	,
(	1580	)	,
(	1583	)	,
(	1587	)	,
(	1590	)	,
(	1594	)	,
(	1597	)	,
(	1601	)	,
(	1604	)	,
(	1608	)	,
(	1611	)	,
(	1615	)	,
(	1618	)	,
(	1622	)	,
(	1625	)	,
(	1629	)	,
(	1632	)	,
(	1636	)	,
(	1639	)	,
(	1642	)	,
(	1646	)	,
(	1649	)	,
(	1653	)	,
(	1656	)	,
(	1660	)	,
(	1663	)	,
(	1666	)	,
(	1670	)	,
(	1673	)	,
(	1677	)	,
(	1680	)	,
(	1683	)	,
(	1687	)	,
(	1690	)	,
(	1693	)	,
(	1697	)	,
(	1700	)	,
(	1704	)	,
(	1707	)	,
(	1710	)	,
(	1714	)	,
(	1717	)	,
(	1720	)	,
(	1723	)	,
(	1727	)	,
(	1730	)	,
(	1733	)	,
(	1737	)	,
(	1740	)	,
(	1743	)	,
(	1747	)	,
(	1750	)	,
(	1753	)	,
(	1756	)	,
(	1760	)	,
(	1763	)	,
(	1766	)	,
(	1769	)	,
(	1773	)	,
(	1776	)	,
(	1779	)	,
(	1782	)	,
(	1786	)	,
(	1789	)	,
(	1792	)	,
(	1795	)	,
(	1798	)	,
(	1802	)	,
(	1805	)	,
(	1808	)	,
(	1811	)	,
(	1814	)	,
(	1817	)	,
(	1821	)	,
(	1824	)	,
(	1827	)	,
(	1830	)	,
(	1833	)	,
(	1836	)	,
(	1840	)	,
(	1843	)	,
(	1846	)	,
(	1849	)	,
(	1852	)	,
(	1855	)	,
(	1858	)	,
(	1861	)	,
(	1864	)	,
(	1868	)	,
(	1871	)	,
(	1874	)	,
(	1877	)	,
(	1880	)	,
(	1883	)	,
(	1886	)	,
(	1889	)	,
(	1892	)	,
(	1895	)	,
(	1898	)	,
(	1901	)	,
(	1904	)	,
(	1907	)	,
(	1910	)	,
(	1914	)	,
(	1917	)	,
(	1920	)	,
(	1923	)	,
(	1926	)	,
(	1929	)	,
(	1932	)	,
(	1935	)	,
(	1938	)	,
(	1941	)	,
(	1944	)	,
(	1947	)	,
(	1950	)	,
(	1953	)	,
(	1956	)	,
(	1958	)	,
(	1961	)	,
(	1964	)	,
(	1967	)	,
(	1970	)	,
(	1973	)	,
(	1976	)	,
(	1979	)	,
(	1982	)	,
(	1985	)	,
(	1988	)	,
(	1991	)	,
(	1994	)	,
(	1997	)	,
(	2000	)	,
(	2003	)	,
(	2005	)	,
(	2008	)	,
(	2011	)	,
(	2014	)	,
(	2017	)	,
(	2020	)	,
(	2023	)	,
(	2026	)	,
(	2029	)	,
(	2031	)	,
(	2034	)	,
(	2037	)	,
(	2040	)	,
(	2043	)	,
(	2046	)	,
(	2049	)	,
(	2051	)	,
(	2054	)	,
(	2057	)	,
(	2060	)	,
(	2063	)	,
(	2065	)	,
(	2068	)	,
(	2071	)	,
(	2074	)	,
(	2077	)	,
(	2080	)	,
(	2082	)	,
(	2085	)	,
(	2088	)	,
(	2091	)	,
(	2094	)	,
(	2096	)	,
(	2099	)	,
(	2102	)	,
(	2105	)	,
(	2107	)	,
(	2110	)	,
(	2113	)	,
(	2116	)	,
(	2118	)	,
(	2121	)	,
(	2124	)	,
(	2127	)	,
(	2129	)	,
(	2132	)	,
(	2135	)	,
(	2138	)	,
(	2140	)	,
(	2143	)	,
(	2146	)	,
(	2148	)	,
(	2151	)	,
(	2154	)	,
(	2157	)	,
(	2159	)	,
(	2162	)	,
(	2165	)	,
(	2167	)	,
(	2170	)	,
(	2173	)	,
(	2175	)	,
(	2178	)	,
(	2181	)	,
(	2183	)	,
(	2186	)	,
(	2189	)	,
(	2191	)	,
(	2194	)	,
(	2197	)	,
(	2199	)	,
(	2202	)	,
(	2205	)	,
(	2207	)	,
(	2210	)	,
(	2213	)	,
(	2215	)	,
(	2218	)	,
(	2220	)	,
(	2223	)	,
(	2226	)	,
(	2228	)	,
(	2231	)	,
(	2234	)	,
(	2236	)	,
(	2239	)	,
(	2241	)	,
(	2244	)	,
(	2247	)	,
(	2249	)	,
(	2252	)	,
(	2254	)	,
(	2257	)	,
(	2259	)	,
(	2262	)	,
(	2265	)	,
(	2267	)	,
(	2270	)	,
(	2272	)	,
(	2275	)	,
(	2277	)	,
(	2280	)	,
(	2282	)	,
(	2285	)	,
(	2288	)	,
(	2290	)	,
(	2293	)	,
(	2295	)	,
(	2298	)	,
(	2300	)	,
(	2303	)	,
(	2305	)	,
(	2308	)	,
(	2310	)	,
(	2313	)	,
(	2315	)	,
(	2318	)	,
(	2320	)	,
(	2323	)	,
(	2325	)	,
(	2328	)	,
(	2330	)	,
(	2333	)	,
(	2335	)	,
(	2338	)	,
(	2340	)	,
(	2343	)	,
(	2345	)	,
(	2348	)	,
(	2350	)	,
(	2353	)	,
(	2355	)	,
(	2357	)	,
(	2360	)	,
(	2362	)	,
(	2365	)	,
(	2367	)	,
(	2370	)	,
(	2372	)	,
(	2375	)	,
(	2377	)	,
(	2379	)	,
(	2382	)	,
(	2384	)	,
(	2387	)	,
(	2389	)	,
(	2392	)	,
(	2394	)	,
(	2396	)	,
(	2399	)	,
(	2401	)	,
(	2404	)	,
(	2406	)	,
(	2408	)	,
(	2411	)	,
(	2413	)	,
(	2416	)	,
(	2418	)	,
(	2420	)	,
(	2423	)	,
(	2425	)	,
(	2428	)	,
(	2430	)	,
(	2432	)	,
(	2435	)	,
(	2437	)	,
(	2439	)	,
(	2442	)	,
(	2444	)	,
(	2447	)	,
(	2449	)	,
(	2451	)	,
(	2454	)	,
(	2456	)	,
(	2458	)	,
(	2461	)	,
(	2463	)	,
(	2465	)	,
(	2468	)	,
(	2470	)	,
(	2472	)	,
(	2475	)	,
(	2477	)	,
(	2479	)	,
(	2482	)	,
(	2484	)	,
(	2486	)	,
(	2489	)	,
(	2491	)	,
(	2493	)	,
(	2495	)	,
(	2498	)	,
(	2500	)	,
(	2502	)	,
(	2505	)	,
(	2507	)	,
(	2509	)	,
(	2511	)	,
(	2514	)	,
(	2516	)	,
(	2518	)	,
(	2521	)	,
(	2523	)	,
(	2525	)	,
(	2527	)	,
(	2530	)	,
(	2532	)	,
(	2534	)	,
(	2536	)	,
(	2539	)	,
(	2541	)	,
(	2543	)	,
(	2545	)	,
(	2548	)	,
(	2550	)	,
(	2552	)	,
(	2554	)	,
(	2557	)	,
(	2559	)	,
(	2561	)	,
(	2563	)	,
(	2566	)	,
(	2568	)	,
(	2570	)	,
(	2572	)	,
(	2575	)	,
(	2577	)	,
(	2579	)	,
(	2581	)	,
(	2583	)	,
(	2586	)	,
(	2588	)	,
(	2590	)	,
(	2592	)	,
(	2594	)	,
(	2597	)	,
(	2599	)	,
(	2601	)	,
(	2603	)	,
(	2605	)	,
(	2608	)	,
(	2610	)	,
(	2612	)	,
(	2614	)	,
(	2616	)	,
(	2618	)	,
(	2621	)	,
(	2623	)	,
(	2625	)	,
(	2627	)	,
(	2629	)	,
(	2631	)	,
(	2634	)	,
(	2636	)	,
(	2638	)	,
(	2640	)	,
(	2642	)	,
(	2644	)	,
(	2647	)	,
(	2649	)	,
(	2651	)	,
(	2653	)	,
(	2655	)	,
(	2657	)	,
(	2659	)	,
(	2661	)	,
(	2664	)	,
(	2666	)	,
(	2668	)	,
(	2670	)	,
(	2672	)	,
(	2674	)	,
(	2676	)	,
(	2678	)	,
(	2681	)	,
(	2683	)	,
(	2685	)	,
(	2687	)	,
(	2689	)	,
(	2691	)	,
(	2693	)	,
(	2695	)	,
(	2697	)	,
(	2699	)	,
(	2702	)	,
(	2704	)	,
(	2706	)	,
(	2708	)	,
(	2710	)	,
(	2712	)	,
(	2714	)	,
(	2716	)	,
(	2718	)	,
(	2720	)	,
(	2722	)	,
(	2724	)	,
(	2726	)	,
(	2729	)	,
(	2731	)	,
(	2733	)	,
(	2735	)	,
(	2737	)	,
(	2739	)	,
(	2741	)	,
(	2743	)	,
(	2745	)	,
(	2747	)	,
(	2749	)	,
(	2751	)	,
(	2753	)	,
(	2755	)	,
(	2757	)	,
(	2759	)	,
(	2761	)	,
(	2763	)	,
(	2765	)	,
(	2767	)	,
(	2769	)	,
(	2771	)	,
(	2773	)	,
(	2775	)	,
(	2777	)	,
(	2779	)	,
(	2782	)	,
(	2784	)	,
(	2786	)	,
(	2788	)	,
(	2790	)	,
(	2792	)	,
(	2794	)	,
(	2796	)	,
(	2798	)	,
(	2800	)	,
(	2802	)	,
(	2804	)	,
(	2806	)	,
(	2808	)	,
(	2809	)	,
(	2811	)	,
(	2813	)	,
(	2815	)	,
(	2817	)	,
(	2819	)	,
(	2821	)	,
(	2823	)	,
(	2825	)	,
(	2827	)	,
(	2829	)	,
(	2831	)	,
(	2833	)	,
(	2835	)	,
(	2837	)	,
(	2839	)	,
(	2841	)	,
(	2843	)	,
(	2845	)	,
(	2847	)	,
(	2849	)	,
(	2851	)	,
(	2853	)	,
(	2855	)	,
(	2857	)	,
(	2859	)	,
(	2861	)	,
(	2862	)	,
(	2864	)	,
(	2866	)	,
(	2868	)	,
(	2870	)	,
(	2872	)	,
(	2874	)	,
(	2876	)	,
(	2878	)	,
(	2880	)	,
(	2882	)	,
(	2884	)	,
(	2886	)	,
(	2887	)	,
(	2889	)	,
(	2891	)	,
(	2893	)	,
(	2895	)	,
(	2897	)	,
(	2899	)	,
(	2901	)	,
(	2903	)	,
(	2905	)	,
(	2907	)	,
(	2908	)	,
(	2910	)	,
(	2912	)	,
(	2914	)	,
(	2916	)	,
(	2918	)	,
(	2920	)	,
(	2922	)	,
(	2924	)	,
(	2925	)	,
(	2927	)	,
(	2929	)	,
(	2931	)	,
(	2933	)	,
(	2935	)	,
(	2937	)	,
(	2939	)	,
(	2940	)	,
(	2942	)	,
(	2944	)	,
(	2946	)	,
(	2948	)	,
(	2950	)	,
(	2952	)	,
(	2953	)	,
(	2955	)	,
(	2957	)	,
(	2959	)	,
(	2961	)	,
(	2963	)	,
(	2965	)	,
(	2966	)	,
(	2968	)	,
(	2970	)	,
(	2972	)	,
(	2974	)	,
(	2976	)	,
(	2977	)	,
(	2979	)	,
(	2981	)	,
(	2983	)	,
(	2985	)	,
(	2987	)	,
(	2988	)	,
(	2990	)	,
(	2992	)	,
(	2994	)	,
(	2996	)	,
(	2997	)	,
(	2999	)	,
(	3001	)	,
(	3003	)	,
(	3005	)	,
(	3007	)	,
(	3008	)	,
(	3010	)	,
(	3012	)	,
(	3014	)	,
(	3016	)	,
(	3017	)	,
(	3019	)	,
(	3021	)	,
(	3023	)	,
(	3025	)	,
(	3026	)	,
(	3028	)	,
(	3030	)	,
(	3032	)	,
(	3034	)	,
(	3035	)	,
(	3037	)	,
(	3039	)	,
(	3041	)	,
(	3042	)	,
(	3044	)	,
(	3046	)	,
(	3048	)	,
(	3050	)	,
(	3051	)	,
(	3053	)	,
(	3055	)	,
(	3057	)	,
(	3058	)	,
(	3060	)	,
(	3062	)	,
(	3064	)	,
(	3065	)	,
(	3067	)	,
(	3069	)	,
(	3071	)	,
(	3072	)	,
(	3074	)	,
(	3076	)	,
(	3078	)	,
(	3079	)	,
(	3081	)	,
(	3083	)	,
(	3085	)	,
(	3086	)	,
(	3088	)	,
(	3090	)	,
(	3092	)	,
(	3093	)	,
(	3095	)	,
(	3097	)	,
(	3099	)	,
(	3100	)	,
(	3102	)	,
(	3104	)	,
(	3106	)	,
(	3107	)	,
(	3109	)	,
(	3111	)	,
(	3112	)	,
(	3114	)	,
(	3116	)	,
(	3118	)	,
(	3119	)	,
(	3121	)	,
(	3123	)	,
(	3124	)	,
(	3126	)	,
(	3128	)	,
(	3130	)	,
(	3131	)	,
(	3133	)	,
(	3135	)	,
(	3136	)	,
(	3138	)	,
(	3140	)	,
(	3142	)	,
(	3143	)	,
(	3145	)	,
(	3147	)	,
(	3148	)	,
(	3150	)	,
(	3152	)	,
(	3153	)	,
(	3155	)	,
(	3157	)	,
(	3158	)	,
(	3160	)	,
(	3162	)	,
(	3163	)	,
(	3165	)	,
(	3167	)	,
(	3169	)	,
(	3170	)	,
(	3172	)	,
(	3174	)	,
(	3175	)	,
(	3177	)	,
(	3179	)	,
(	3180	)	,
(	3182	)	,
(	3184	)	,
(	3185	)	,
(	3187	)	,
(	3189	)	,
(	3190	)	,
(	3192	)	,
(	3194	)	,
(	3195	)	,
(	3197	)	,
(	3198	)	,
(	3200	)	,
(	3202	)	,
(	3203	)	,
(	3205	)	,
(	3207	)	,
(	3208	)	,
(	3210	)	,
(	3212	)	,
(	3213	)	,
(	3215	)	,
(	3217	)	,
(	3218	)	,
(	3220	)	,
(	3221	)	,
(	3223	)	,
(	3225	)	,
(	3226	)	,
(	3228	)	,
(	3230	)	,
(	3231	)	,
(	3233	)	,
(	3235	)	,
(	3236	)	,
(	3238	)	,
(	3239	)	,
(	3241	)	,
(	3243	)	,
(	3244	)	,
(	3246	)	,
(	3247	)	,
(	3249	)	,
(	3251	)	,
(	3252	)	,
(	3254	)	,
(	3256	)	,
(	3257	)	,
(	3259	)	,
(	3260	)	,
(	3262	)	,
(	3264	)	,
(	3265	)	,
(	3267	)	,
(	3268	)	,
(	3270	)	,
(	3272	)	,
(	3273	)	,
(	3275	)	,
(	3276	)	,
(	3278	)	,
(	3280	)	,
(	3281	)	,
(	3283	)	,
(	3284	)	,
(	3286	)	,
(	3287	)	,
(	3289	)	,
(	3291	)	,
(	3292	)	,
(	3294	)	,
(	3295	)	,
(	3297	)	,
(	3299	)	,
(	3300	)	,
(	3302	)	,
(	3303	)	,
(	3305	)	,
(	3306	)	,
(	3308	)	,
(	3310	)	,
(	3311	)	,
(	3313	)	,
(	3314	)	,
(	3316	)	,
(	3317	)	,
(	3319	)	,
(	3321	)	,
(	3322	)	,
(	3324	)	,
(	3325	)	,
(	3327	)	,
(	3328	)	,
(	3330	)	,
(	3331	)	,
(	3333	)	,
(	3335	)	,
(	3336	)	,
(	3338	)	,
(	3339	)	,
(	3341	)	,
(	3342	)	,
(	3344	)	,
(	3345	)	,
(	3347	)	,
(	3348	)	,
(	3350	)	,
(	3352	)	,
(	3353	)	,
(	3355	)	,
(	3356	)	,
(	3358	)	,
(	3359	)	,
(	3361	)	,
(	3362	)	,
(	3364	)	,
(	3365	)	,
(	3367	)	,
(	3368	)	,
(	3370	)	,
(	3371	)	,
(	3373	)	,
(	3374	)	,
(	3376	)	,
(	3377	)	,
(	3379	)	,
(	3381	)	,
(	3382	)	,
(	3384	)	,
(	3385	)	,
(	3387	)	,
(	3388	)	,
(	3390	)	,
(	3391	)	,
(	3393	)	,
(	3394	)	,
(	3396	)	,
(	3397	)	,
(	3399	)	,
(	3400	)	,
(	3402	)	,
(	3403	)	,
(	3405	)	,
(	3406	)	,
(	3408	)	,
(	3409	)	,
(	3411	)	,
(	3412	)	,
(	3414	)	,
(	3415	)	,
(	3417	)	,
(	3418	)	,
(	3420	)	,
(	3421	)	,
(	3423	)	,
(	3424	)	,
(	3426	)	,
(	3427	)	,
(	3429	)	,
(	3430	)	,
(	3431	)	,
(	3433	)	,
(	3434	)	,
(	3436	)	,
(	3437	)	,
(	3439	)	,
(	3440	)	,
(	3442	)	,
(	3443	)	,
(	3445	)	,
(	3446	)	,
(	3448	)	,
(	3449	)	,
(	3451	)	,
(	3452	)	,
(	3454	)	,
(	3455	)	,
(	3457	)	,
(	3458	)	,
(	3459	)	,
(	3461	)	,
(	3462	)	,
(	3464	)	,
(	3465	)	,
(	3467	)	,
(	3468	)	,
(	3470	)	,
(	3471	)	,
(	3473	)	,
(	3474	)	,
(	3475	)	,
(	3477	)	,
(	3478	)	,
(	3480	)	,
(	3481	)	,
(	3483	)	,
(	3484	)	,
(	3486	)	,
(	3487	)	,
(	3488	)	,
(	3490	)	,
(	3491	)	,
(	3493	)	,
(	3494	)	,
(	3496	)	,
(	3497	)	,
(	3499	)	,
(	3500	)	,
(	3501	)	,
(	3503	)	,
(	3504	)	,
(	3506	)	,
(	3507	)	,
(	3509	)	,
(	3510	)	,
(	3511	)	,
(	3513	)	,
(	3514	)	,
(	3516	)	,
(	3517	)	,
(	3519	)	,
(	3520	)	,
(	3521	)	,
(	3523	)	,
(	3524	)	,
(	3526	)	,
(	3527	)	,
(	3528	)	,
(	3530	)	,
(	3531	)	,
(	3533	)	,
(	3534	)	,
(	3536	)	,
(	3537	)	,
(	3538	)	,
(	3540	)	,
(	3541	)	,
(	3543	)	,
(	3544	)	,
(	3545	)	,
(	3547	)	,
(	3548	)	,
(	3550	)	,
(	3551	)	,
(	3552	)	,
(	3554	)	,
(	3555	)	,
(	3557	)	,
(	3558	)	,
(	3559	)	,
(	3561	)	,
(	3562	)	,
(	3564	)	,
(	3565	)	,
(	3566	)	,
(	3568	)	,
(	3569	)	,
(	3570	)	,
(	3572	)	,
(	3573	)	,
(	3575	)	,
(	3576	)	,
(	3577	)	,
(	3579	)	,
(	3580	)	,
(	3582	)	,
(	3583	)	,
(	3584	)	,
(	3586	)	,
(	3587	)	,
(	3588	)	,
(	3590	)	,
(	3591	)	,
(	3593	)	,
(	3594	)	,
(	3595	)	,
(	3597	)	,
(	3598	)	,
(	3599	)	,
(	3601	)	,
(	3602	)	,
(	3604	)	,
(	3605	)	,
(	3606	)	,
(	3608	)	,
(	3609	)	,
(	3610	)	,
(	3612	)	,
(	3613	)	,
(	3614	)	,
(	3616	)	,
(	3617	)	,
(	3618	)	,
(	3620	)	,
(	3621	)	,
(	3623	)	,
(	3624	)	,
(	3625	)	,
(	3627	)	,
(	3628	)	,
(	3629	)	,
(	3631	)	,
(	3632	)	,
(	3633	)	,
(	3635	)	,
(	3636	)	,
(	3637	)	,
(	3639	)	,
(	3640	)	,
(	3641	)	,
(	3643	)	,
(	3644	)	,
(	3645	)	,
(	3647	)	,
(	3648	)	,
(	3649	)	,
(	3651	)	,
(	3652	)	,
(	3653	)	,
(	3655	)	,
(	3656	)	,
(	3657	)	,
(	3659	)	,
(	3660	)	,
(	3661	)	,
(	3663	)	,
(	3664	)	,
(	3665	)	,
(	3667	)	,
(	3668	)	,
(	3669	)	,
(	3671	)	,
(	3672	)	,
(	3673	)	,
(	3675	)	,
(	3676	)	,
(	3677	)	,
(	3679	)	,
(	3680	)	,
(	3681	)	,
(	3683	)	,
(	3684	)	,
(	3685	)	,
(	3687	)	,
(	3688	)	,
(	3689	)	,
(	3690	)	,
(	3692	)	,
(	3693	)	,
(	3694	)	,
(	3696	)	,
(	3697	)	,
(	3698	)	,
(	3700	)	,
(	3701	)	,
(	3702	)	,
(	3704	)	,
(	3705	)	,
(	3706	)	,
(	3707	)	,
(	3709	)	,
(	3710	)	,
(	3711	)	,
(	3713	)	,
(	3714	)	,
(	3715	)	,
(	3717	)	,
(	3718	)	,
(	3719	)	,
(	3720	)	,
(	3722	)	,
(	3723	)	,
(	3724	)	,
(	3726	)	,
(	3727	)	,
(	3728	)	,
(	3729	)	,
(	3731	)	,
(	3732	)	,
(	3733	)	,
(	3735	)	,
(	3736	)	,
(	3737	)	,
(	3738	)	,
(	3740	)	,
(	3741	)	,
(	3742	)	,
(	3744	)	,
(	3745	)	,
(	3746	)	,
(	3747	)	,
(	3749	)	,
(	3750	)	,
(	3751	)	,
(	3752	)	,
(	3754	)	,
(	3755	)	,
(	3756	)	,
(	3758	)	,
(	3759	)	,
(	3760	)	,
(	3761	)	,
(	3763	)	,
(	3764	)	,
(	3765	)	,
(	3766	)	,
(	3768	)	,
(	3769	)	,
(	3770	)	,
(	3771	)	,
(	3773	)	,
(	3774	)	,
(	3775	)	,
(	3777	)	,
(	3778	)	,
(	3779	)	,
(	3780	)	,
(	3782	)	,
(	3783	)	,
(	3784	)	,
(	3785	)	,
(	3787	)	,
(	3788	)	,
(	3789	)	,
(	3790	)	,
(	3792	)	,
(	3793	)	,
(	3794	)	,
(	3795	)	,
(	3797	)	,
(	3798	)	,
(	3799	)	,
(	3800	)	,
(	3802	)	,
(	3803	)	,
(	3804	)	,
(	3805	)	,
(	3807	)	,
(	3808	)	,
(	3809	)	,
(	3810	)	,
(	3811	)	,
(	3813	)	,
(	3814	)	,
(	3815	)	,
(	3816	)	,
(	3818	)	,
(	3819	)	,
(	3820	)	,
(	3821	)	,
(	3823	)	,
(	3824	)	,
(	3825	)	,
(	3826	)	,
(	3828	)	,
(	3829	)	,
(	3830	)	,
(	3831	)	,
(	3832	)	,
(	3834	)	,
(	3835	)	,
(	3836	)	,
(	3837	)	,
(	3839	)	,
(	3840	)	,
(	3841	)	,
(	3842	)	,
(	3843	)	,
(	3845	)	,
(	3846	)	,
(	3847	)	,
(	3848	)	,
(	3850	)	,
(	3851	)	,
(	3852	)	,
(	3853	)	,
(	3854	)	,
(	3856	)	,
(	3857	)	,
(	3858	)	,
(	3859	)	,
(	3860	)	,
(	3862	)	,
(	3863	)	,
(	3864	)	,
(	3865	)	,
(	3866	)	,
(	3868	)	,
(	3869	)	,
(	3870	)	,
(	3871	)	,
(	3872	)	,
(	3874	)	,
(	3875	)	,
(	3876	)	,
(	3877	)	,
(	3879	)	,
(	3880	)	,
(	3881	)	,
(	3882	)	,
(	3883	)	,
(	3884	)	,
(	3886	)	,
(	3887	)	,
(	3888	)	,
(	3889	)	,
(	3890	)	,
(	3892	)	,
(	3893	)	,
(	3894	)	,
(	3895	)	,
(	3896	)	,
(	3898	)	,
(	3899	)	,
(	3900	)	,
(	3901	)	,
(	3902	)	,
(	3904	)	,
(	3905	)	,
(	3906	)	,
(	3907	)	,
(	3908	)	,
(	3909	)	,
(	3911	)	,
(	3912	)	,
(	3913	)	,
(	3914	)	,
(	3915	)	,
(	3917	)	,
(	3918	)	,
(	3919	)	,
(	3920	)	,
(	3921	)	,
(	3922	)	,
(	3924	)	,
(	3925	)	,
(	3926	)	,
(	3927	)	,
(	3928	)	,
(	3929	)	,
(	3931	)	,
(	3932	)	,
(	3933	)	,
(	3934	)	,
(	3935	)	,
(	3936	)	,
(	3938	)	,
(	3939	)	,
(	3940	)	,
(	3941	)	,
(	3942	)	,
(	3943	)	,
(	3945	)	,
(	3946	)	,
(	3947	)	,
(	3948	)	,
(	3949	)	,
(	3950	)	,
(	3952	)	,
(	3953	)	,
(	3954	)	,
(	3955	)	,
(	3956	)	,
(	3957	)	,
(	3959	)	,
(	3960	)	,
(	3961	)	,
(	3962	)	,
(	3963	)	,
(	3964	)	,
(	3965	)	,
(	3967	)	,
(	3968	)	,
(	3969	)	,
(	3970	)	,
(	3971	)	,
(	3972	)	,
(	3974	)	,
(	3975	)	,
(	3976	)	,
(	3977	)	,
(	3978	)	,
(	3979	)	,
(	3980	)	,
(	3982	)	,
(	3983	)	,
(	3984	)	,
(	3985	)	,
(	3986	)	,
(	3987	)	,
(	3988	)	,
(	3990	)	,
(	3991	)	,
(	3992	)	,
(	3993	)	,
(	3994	)	,
(	3995	)	,
(	3996	)	,
(	3997	)	,
(	3999	)	,
(	4000	)	,
(	4001	)	,
(	4002	)	,
(	4003	)	,
(	4004	)	,
(	4005	)	,
(	4007	)	,
(	4008	)	,
(	4009	)	,
(	4010	)	,
(	4011	)	,
(	4012	)	,
(	4013	)	,
(	4014	)	,
(	4016	)	,
(	4017	)	,
(	4018	)	,
(	4019	)	,
(	4020	)	,
(	4021	)	,
(	4022	)	,
(	4023	)	,
(	4025	)	,
(	4026	)	,
(	4027	)	,
(	4028	)	,
(	4029	)	,
(	4030	)	,
(	4031	)	,
(	4032	)	,
(	4033	)	,
(	4035	)	,
(	4036	)	,
(	4037	)	,
(	4038	)	,
(	4039	)	,
(	4040	)	,
(	4041	)	,
(	4042	)	,
(	4043	)	,
(	4045	)	,
(	4046	)	,
(	4047	)	,
(	4048	)	,
(	4049	)	,
(	4050	)	,
(	4051	)	,
(	4052	)	,
(	4053	)	,
(	4055	)	,
(	4056	)	,
(	4057	)	,
(	4058	)	,
(	4059	)	,
(	4060	)	,
(	4061	)	,
(	4062	)	,
(	4063	)	,
(	4064	)	,
(	4066	)	,
(	4067	)	,
(	4068	)	,
(	4069	)	,
(	4070	)	,
(	4071	)	,
(	4072	)	,
(	4073	)	,
(	4074	)	,
(	4075	)	,
(	4076	)	,
(	4078	)	,
(	4079	)	,
(	4080	)	,
(	4081	)	,
(	4082	)	,
(	4083	)	,
(	4084	)	,
(	4085	)	,
(	4086	)	,
(	4087	)	,
(	4088	)	,
(	4090	)	,
(	4091	)	,
(	4092	)	,
(	4093	)	,
(	4094	)	,
(	4095	)	,
(	4096	)	,
(	4097	)	,
(	4098	)	,
(	4099	)	,
(	4100	)	,
(	4101	)	,
(	4103	)	,
(	4104	)	,
(	4105	)	,
(	4106	)	,
(	4107	)	,
(	4108	)	,
(	4109	)	,
(	4110	)	,
(	4111	)	,
(	4112	)	,
(	4113	)	,
(	4114	)	,
(	4115	)	,
(	4117	)	,
(	4118	)	,
(	4119	)	,
(	4120	)	,
(	4121	)	,
(	4122	)	,
(	4123	)	,
(	4124	)	,
(	4125	)	,
(	4126	)	,
(	4127	)	,
(	4128	)	,
(	4129	)	,
(	4130	)	,
(	4131	)	,
(	4133	)	,
(	4134	)	,
(	4135	)	,
(	4136	)	,
(	4137	)	,
(	4138	)	,
(	4139	)	,
(	4140	)	,
(	4141	)	,
(	4142	)	,
(	4143	)	,
(	4144	)	,
(	4145	)	,
(	4146	)	,
(	4147	)	,
(	4148	)	,
(	4150	)	,
(	4151	)	,
(	4152	)	,
(	4153	)	,
(	4154	)	,
(	4155	)	,
(	4156	)	,
(	4157	)	,
(	4158	)	,
(	4159	)	,
(	4160	)	,
(	4161	)	,
(	4162	)	,
(	4163	)	,
(	4164	)	,
(	4165	)	,
(	4166	)	,
(	4167	)	,
(	4168	)	,
(	4169	)	,
(	4171	)	,
(	4172	)	,
(	4173	)	,
(	4174	)	,
(	4175	)	,
(	4176	)	,
(	4177	)	,
(	4178	)	,
(	4179	)	,
(	4180	)	,
(	4181	)	,
(	4182	)	,
(	4183	)	,
(	4184	)	,
(	4185	)	,
(	4186	)	,
(	4187	)	,
(	4188	)	,
(	4189	)	,
(	4190	)	,
(	4191	)	,
(	4192	)	,
(	4193	)	,
(	4194	)	,
(	4195	)	,
(	4196	)	,
(	4198	)	,
(	4199	)	,
(	4200	)	,
(	4201	)	,
(	4202	)	,
(	4203	)	,
(	4204	)	,
(	4205	)	,
(	4206	)	,
(	4207	)	,
(	4208	)	,
(	4209	)	,
(	4210	)	,
(	4211	)	,
(	4212	)	,
(	4213	)	,
(	4214	)	,
(	4215	)	,
(	4216	)	,
(	4217	)	,
(	4218	)	,
(	4219	)	,
(	4220	)	,
(	4221	)	,
(	4222	)	,
(	4223	)	,
(	4224	)	,
(	4225	)	,
(	4226	)	,
(	4227	)	,
(	4228	)	,
(	4229	)	,
(	4230	)	,
(	4231	)	,
(	4232	)	,
(	4233	)	,
(	4234	)	,
(	4235	)	,
(	4236	)	,
(	4237	)	,
(	4238	)	,
(	4239	)	,
(	4240	)	,
(	4241	)	,
(	4242	)	,
(	4243	)	,
(	4244	)	,
(	4245	)	,
(	4246	)	,
(	4248	)	,
(	4249	)	,
(	4250	)	,
(	4251	)	,
(	4252	)	,
(	4253	)	,
(	4254	)	,
(	4255	)	,
(	4256	)	,
(	4257	)	,
(	4258	)	,
(	4259	)	,
(	4260	)	,
(	4261	)	,
(	4262	)	,
(	4263	)	,
(	4264	)	,
(	4265	)	,
(	4266	)	,
(	4267	)	,
(	4268	)	,
(	4269	)	,
(	4270	)	,
(	4271	)	,
(	4272	)	,
(	4273	)	,
(	4274	)	,
(	4275	)	,
(	4276	)	,
(	4277	)	,
(	4278	)	,
(	4279	)	,
(	4280	)	,
(	4281	)	,
(	4282	)	,
(	4282	)	,
(	4283	)	,
(	4284	)	,
(	4285	)	,
(	4286	)	,
(	4287	)	,
(	4288	)	,
(	4289	)	,
(	4290	)	,
(	4291	)	,
(	4292	)	,
(	4293	)	,
(	4294	)	,
(	4295	)	,
(	4296	)	,
(	4297	)	,
(	4298	)	,
(	4299	)	,
(	4300	)	,
(	4301	)	,
(	4302	)	,
(	4303	)	,
(	4304	)	,
(	4305	)	,
(	4306	)	,
(	4307	)	,
(	4308	)	,
(	4309	)	,
(	4310	)	,
(	4311	)	,
(	4312	)	,
(	4313	)	,
(	4314	)	,
(	4315	)	,
(	4316	)	,
(	4317	)	,
(	4318	)	,
(	4319	)	,
(	4320	)	,
(	4321	)	,
(	4322	)	,
(	4323	)	,
(	4324	)	,
(	4325	)	,
(	4326	)	,
(	4327	)	,
(	4328	)	,
(	4329	)	,
(	4330	)	,
(	4331	)	,
(	4331	)	,
(	4332	)	,
(	4333	)	,
(	4334	)	,
(	4335	)	,
(	4336	)	,
(	4337	)	,
(	4338	)	,
(	4339	)	,
(	4340	)	,
(	4341	)	,
(	4342	)	,
(	4343	)	,
(	4344	)	,
(	4345	)	,
(	4346	)	,
(	4347	)	,
(	4348	)	,
(	4349	)	,
(	4350	)	,
(	4351	)	,
(	4352	)	,
(	4353	)	,
(	4354	)	,
(	4355	)	,
(	4356	)	,
(	4357	)	,
(	4357	)	,
(	4358	)	,
(	4359	)	,
(	4360	)	,
(	4361	)	,
(	4362	)	,
(	4363	)	,
(	4364	)	,
(	4365	)	,
(	4366	)	,
(	4367	)	,
(	4368	)	,
(	4369	)	,
(	4370	)	,
(	4371	)	,
(	4372	)	,
(	4373	)	,
(	4374	)	,
(	4375	)	,
(	4376	)	,
(	4377	)	,
(	4377	)	,
(	4378	)	,
(	4379	)	,
(	4380	)	,
(	4381	)	,
(	4382	)	,
(	4383	)	,
(	4384	)	,
(	4385	)	,
(	4386	)	,
(	4387	)	,
(	4388	)	,
(	4389	)	,
(	4390	)	,
(	4391	)	,
(	4392	)	,
(	4393	)	,
(	4394	)	,
(	4394	)	,
(	4395	)	,
(	4396	)	,
(	4397	)	,
(	4398	)	,
(	4399	)	,
(	4400	)	,
(	4401	)	,
(	4402	)	,
(	4403	)	,
(	4404	)	,
(	4405	)	,
(	4406	)	,
(	4407	)	,
(	4408	)	,
(	4409	)	,
(	4409	)	,
(	4410	)	,
(	4411	)	,
(	4412	)	,
(	4413	)	,
(	4414	)	,
(	4415	)	,
(	4416	)	,
(	4417	)	,
(	4418	)	,
(	4419	)	,
(	4420	)	,
(	4421	)	,
(	4422	)	,
(	4423	)	,
(	4423	)	,
(	4424	)	,
(	4425	)	,
(	4426	)	,
(	4427	)	,
(	4428	)	,
(	4429	)	,
(	4430	)	,
(	4431	)	,
(	4432	)	,
(	4433	)	,
(	4434	)	,
(	4435	)	,
(	4435	)	,
(	4436	)	,
(	4437	)	,
(	4438	)	,
(	4439	)	,
(	4440	)	,
(	4441	)	,
(	4442	)	,
(	4443	)	,
(	4444	)	,
(	4445	)	,
(	4446	)	,
(	4447	)	,
(	4447	)	,
(	4448	)	,
(	4449	)	,
(	4450	)	,
(	4451	)	,
(	4452	)	,
(	4453	)	,
(	4454	)	,
(	4455	)	,
(	4456	)	,
(	4457	)	,
(	4458	)	,
(	4458	)	,
(	4459	)	,
(	4460	)	,
(	4461	)	,
(	4462	)	,
(	4463	)	,
(	4464	)	,
(	4465	)	,
(	4466	)	,
(	4467	)	,
(	4468	)	,
(	4468	)	,
(	4469	)	,
(	4470	)	,
(	4471	)	,
(	4472	)	,
(	4473	)	,
(	4474	)	,
(	4475	)	,
(	4476	)	,
(	4477	)	,
(	4477	)	,
(	4478	)	,
(	4479	)	,
(	4480	)	,
(	4481	)	,
(	4482	)	,
(	4483	)	,
(	4484	)	,
(	4485	)	,
(	4486	)	,
(	4487	)	,
(	4487	)	,
(	4488	)	,
(	4489	)	,
(	4490	)	,
(	4491	)	,
(	4492	)	,
(	4493	)	,
(	4494	)	,
(	4495	)	,
(	4496	)	,
(	4496	)	,
(	4497	)	,
(	4498	)	,
(	4499	)	,
(	4500	)	,
(	4501	)	,
(	4502	)	,
(	4503	)	,
(	4504	)	,
(	4504	)	,
(	4505	)	,
(	4506	)	,
(	4507	)	,
(	4508	)	,
(	4509	)	,
(	4510	)	,
(	4511	)	,
(	4512	)	,
(	4512	)	,
(	4513	)	,
(	4514	)	,
(	4515	)	,
(	4516	)	,
(	4517	)	,
(	4518	)	,
(	4519	)	,
(	4520	)	,
(	4520	)	,
(	4521	)	,
(	4522	)	,
(	4523	)	,
(	4524	)	,
(	4525	)	,
(	4526	)	,
(	4527	)	,
(	4528	)	,
(	4528	)	,
(	4529	)	,
(	4530	)	,
(	4531	)	,
(	4532	)	,
(	4533	)	,
(	4534	)	,
(	4535	)	,
(	4535	)	,
(	4536	)	,
(	4537	)	,
(	4538	)	,
(	4539	)	,
(	4540	)	,
(	4541	)	,
(	4542	)	,
(	4543	)	,
(	4543	)	,
(	4544	)	,
(	4545	)	,
(	4546	)	,
(	4547	)	,
(	4548	)	,
(	4549	)	,
(	4550	)	,
(	4550	)	,
(	4551	)	,
(	4552	)	,
(	4553	)	,
(	4554	)	,
(	4555	)	,
(	4556	)	,
(	4556	)	,
(	4557	)	,
(	4558	)	,
(	4559	)	,
(	4560	)	,
(	4561	)	,
(	4562	)	,
(	4563	)	,
(	4563	)	,
(	4564	)	,
(	4565	)	,
(	4566	)	,
(	4567	)	,
(	4568	)	,
(	4569	)	,
(	4570	)	,
(	4570	)	,
(	4571	)	,
(	4572	)	,
(	4573	)	,
(	4574	)	,
(	4575	)	,
(	4576	)	,
(	4576	)	,
(	4577	)	,
(	4578	)	,
(	4579	)	,
(	4580	)	,
(	4581	)	,
(	4582	)	,
(	4582	)	,
(	4583	)	,
(	4584	)	,
(	4585	)	,
(	4586	)	,
(	4587	)	,
(	4588	)	,
(	4588	)	,
(	4589	)	,
(	4590	)	,
(	4591	)	,
(	4592	)	,
(	4593	)	,
(	4594	)	,
(	4594	)	,
(	4595	)	,
(	4596	)	,
(	4597	)	,
(	4598	)	,
(	4599	)	,
(	4600	)	,
(	4600	)	,
(	4601	)	,
(	4602	)	,
(	4603	)	,
(	4604	)	,
(	4605	)	,
(	4606	)	,
(	4606	)	,
(	4607	)	,
(	4608	)	,
(	4609	)	,
(	4610	)	,
(	4611	)	,
(	4612	)	,
(	4612	)	,
(	4613	)	,
(	4614	)	,
(	4615	)	,
(	4616	)	,
(	4617	)	,
(	4617	)	,
(	4618	)	,
(	4619	)	,
(	4620	)	,
(	4621	)	,
(	4622	)	,
(	4623	)	,
(	4623	)	,
(	4624	)	,
(	4625	)	,
(	4626	)	,
(	4627	)	,
(	4628	)	,
(	4628	)	,
(	4629	)	,
(	4630	)	,
(	4631	)	,
(	4632	)	,
(	4633	)	,
(	4633	)	,
(	4634	)	,
(	4635	)	,
(	4636	)	,
(	4637	)	,
(	4638	)	,
(	4639	)	,
(	4639	)	,
(	4640	)	,
(	4641	)	,
(	4642	)	,
(	4643	)	,
(	4644	)	,
(	4644	)	,
(	4645	)	,
(	4646	)	,
(	4647	)	,
(	4648	)	,
(	4649	)	,
(	4649	)	,
(	4650	)	,
(	4651	)	,
(	4652	)	,
(	4653	)	,
(	4654	)	,
(	4654	)	,
(	4655	)	,
(	4656	)	,
(	4657	)	,
(	4658	)	,
(	4659	)	,
(	4659	)	,
(	4660	)	,
(	4661	)	,
(	4662	)	,
(	4663	)	,
(	4664	)	,
(	4664	)	,
(	4665	)	,
(	4666	)	,
(	4667	)	,
(	4668	)	,
(	4668	)	,
(	4669	)	,
(	4670	)	,
(	4671	)	,
(	4672	)	,
(	4673	)	,
(	4673	)	,
(	4674	)	,
(	4675	)	,
(	4676	)	,
(	4677	)	,
(	4678	)	,
(	4678	)	,
(	4679	)	,
(	4680	)	,
(	4681	)	,
(	4682	)	,
(	4683	)	,
(	4683	)	,
(	4684	)	,
(	4685	)	,
(	4686	)	,
(	4687	)	,
(	4687	)	,
(	4688	)	,
(	4689	)	,
(	4690	)	,
(	4691	)	,
(	4692	)	,
(	4692	)	,
(	4693	)	,
(	4694	)	,
(	4695	)	,
(	4696	)	,
(	4696	)	,
(	4697	)	,
(	4698	)	,
(	4699	)	,
(	4700	)	,
(	4700	)	,
(	4701	)	,
(	4702	)	,
(	4703	)	,
(	4704	)	,
(	4705	)	,
(	4705	)	,
(	4706	)	,
(	4707	)	,
(	4708	)	,
(	4709	)	,
(	4709	)	,
(	4710	)	,
(	4711	)	,
(	4712	)	,
(	4713	)	,
(	4713	)	,
(	4714	)	,
(	4715	)	,
(	4716	)	,
(	4717	)	,
(	4718	)	,
(	4718	)	,
(	4719	)	,
(	4720	)	,
(	4721	)	,
(	4722	)	,
(	4722	)	,
(	4723	)	,
(	4724	)	,
(	4725	)	,
(	4726	)	,
(	4726	)	,
(	4727	)	,
(	4728	)	,
(	4729	)	,
(	4730	)	,
(	4730	)	,
(	4731	)	,
(	4732	)	,
(	4733	)	,
(	4734	)	,
(	4734	)	,
(	4735	)	,
(	4736	)	,
(	4737	)	,
(	4738	)	,
(	4738	)	,
(	4739	)	,
(	4740	)	,
(	4741	)	,
(	4742	)	,
(	4742	)	,
(	4743	)	,
(	4744	)	,
(	4745	)	,
(	4746	)	,
(	4746	)	,
(	4747	)	,
(	4748	)	,
(	4749	)	,
(	4750	)	,
(	4750	)	,
(	4751	)	,
(	4752	)	,
(	4753	)	,
(	4754	)	,
(	4754	)	,
(	4755	)	,
(	4756	)	,
(	4757	)	,
(	4758	)	,
(	4758	)	,
(	4759	)	,
(	4760	)	,
(	4761	)	,
(	4761	)	,
(	4762	)	,
(	4763	)	,
(	4764	)	,
(	4765	)	,
(	4765	)	,
(	4766	)	,
(	4767	)	,
(	4768	)	,
(	4769	)	,
(	4769	)	,
(	4770	)	,
(	4771	)	,
(	4772	)	,
(	4773	)	,
(	4773	)	,
(	4774	)	,
(	4775	)	,
(	4776	)	,
(	4776	)	,
(	4777	)	,
(	4778	)	,
(	4779	)	,
(	4780	)	,
(	4780	)	,
(	4781	)	,
(	4782	)	,
(	4783	)	,
(	4784	)	,
(	4784	)	,
(	4785	)	,
(	4786	)	,
(	4787	)	,
(	4787	)	,
(	4788	)	,
(	4789	)	,
(	4790	)	,
(	4791	)	,
(	4791	)	,
(	4792	)	,
(	4793	)	,
(	4794	)	,
(	4794	)	,
(	4795	)	,
(	4796	)	,
(	4797	)	,
(	4798	)	,
(	4798	)	,
(	4799	)	,
(	4800	)	,
(	4801	)	,
(	4801	)	,
(	4802	)	,
(	4803	)	,
(	4804	)	,
(	4805	)	,
(	4805	)	,
(	4806	)	,
(	4807	)	,
(	4808	)	,
(	4808	)	,
(	4809	)	,
(	4810	)	,
(	4811	)	,
(	4812	)	,
(	4812	)	,
(	4813	)	,
(	4814	)	,
(	4815	)	,
(	4815	)	,
(	4816	)	,
(	4817	)	,
(	4818	)	,
(	4818	)	,
(	4819	)	,
(	4820	)	,
(	4821	)	,
(	4822	)	,
(	4822	)	,
(	4823	)	,
(	4824	)	,
(	4825	)	,
(	4825	)	,
(	4826	)	,
(	4827	)	,
(	4828	)	,
(	4828	)	,
(	4829	)	,
(	4830	)	,
(	4831	)	,
(	4832	)	,
(	4832	)	,
(	4833	)	,
(	4834	)	,
(	4835	)	,
(	4835	)	,
(	4836	)	,
(	4837	)	,
(	4838	)	,
(	4838	)	,
(	4839	)	,
(	4840	)	,
(	4841	)	,
(	4841	)	,
(	4842	)	,
(	4843	)	,
(	4844	)	,
(	4844	)	,
(	4845	)	,
(	4846	)	,
(	4847	)	,
(	4848	)	,
(	4848	)	,
(	4849	)	,
(	4850	)	,
(	4851	)	,
(	4851	)	,
(	4852	)	,
(	4853	)	,
(	4854	)	,
(	4854	)	,
(	4855	)	,
(	4856	)	,
(	4857	)	,
(	4857	)	,
(	4858	)	,
(	4859	)	,
(	4860	)	,
(	4860	)	,
(	4861	)	,
(	4862	)	,
(	4863	)	,
(	4863	)	,
(	4864	)	,
(	4865	)	,
(	4866	)	,
(	4866	)	,
(	4867	)	,
(	4868	)	,
(	4869	)	,
(	4869	)	,
(	4870	)	,
(	4871	)	,
(	4872	)	,
(	4872	)	,
(	4873	)	,
(	4874	)	,
(	4875	)	,
(	4875	)	,
(	4876	)	,
(	4877	)	,
(	4878	)	,
(	4878	)	,
(	4879	)	,
(	4880	)	,
(	4881	)	,
(	4881	)	,
(	4882	)	,
(	4883	)	,
(	4884	)	,
(	4884	)	,
(	4885	)	,
(	4886	)	,
(	4887	)	,
(	4887	)	,
(	4888	)	,
(	4889	)	,
(	4890	)	,
(	4890	)	,
(	4891	)	,
(	4892	)	,
(	4893	)	,
(	4893	)	,
(	4894	)	,
(	4895	)	,
(	4896	)	,
(	4896	)	,
(	4897	)	,
(	4898	)	,
(	4899	)	,
(	4899	)	,
(	4900	)	,
(	4901	)	,
(	4902	)	,
(	4902	)	,
(	4903	)	,
(	4904	)	,
(	4904	)	,
(	4905	)	,
(	4906	)	,
(	4907	)	,
(	4907	)	,
(	4908	)	,
(	4909	)	,
(	4910	)	,
(	4910	)	,
(	4911	)	,
(	4912	)	,
(	4913	)	,
(	4913	)	,
(	4914	)	,
(	4915	)	,
(	4916	)	,
(	4916	)	,
(	4917	)	,
(	4918	)	,
(	4918	)	,
(	4919	)	,
(	4920	)	,
(	4921	)	,
(	4921	)	,
(	4922	)	,
(	4923	)	,
(	4924	)	,
(	4924	)	,
(	4925	)	,
(	4926	)	,
(	4927	)	,
(	4927	)	,
(	4928	)	,
(	4929	)	,
(	4929	)	,
(	4930	)	,
(	4931	)	,
(	4932	)	,
(	4932	)	,
(	4933	)	,
(	4934	)	,
(	4935	)	,
(	4935	)	,
(	4936	)	,
(	4937	)	,
(	4937	)	,
(	4938	)	,
(	4939	)	,
(	4940	)	,
(	4940	)	,
(	4941	)	,
(	4942	)	,
(	4943	)	,
(	4943	)	,
(	4944	)	,
(	4945	)	,
(	4945	)	,
(	4946	)	,
(	4947	)	,
(	4948	)	,
(	4948	)	,
(	4949	)	,
(	4950	)	,
(	4951	)	,
(	4951	)	,
(	4952	)	,
(	4953	)	,
(	4953	)	,
(	4954	)	,
(	4955	)	,
(	4956	)	,
(	4956	)	,
(	4957	)	,
(	4958	)	,
(	4959	)	,
(	4959	)	,
(	4960	)	,
(	4961	)	,
(	4961	)	,
(	4962	)	,
(	4963	)	,
(	4964	)	,
(	4964	)	,
(	4965	)	,
(	4966	)	,
(	4966	)	,
(	4967	)	,
(	4968	)	,
(	4969	)	,
(	4969	)	,
(	4970	)	,
(	4971	)	,
(	4971	)	,
(	4972	)	,
(	4973	)	,
(	4974	)	,
(	4974	)	,
(	4975	)	,
(	4976	)	,
(	4976	)	,
(	4977	)	,
(	4978	)	,
(	4979	)	,
(	4979	)	,
(	4980	)	,
(	4981	)	,
(	4981	)	,
(	4982	)	,
(	4983	)	,
(	4984	)	,
(	4984	)	,
(	4985	)	,
(	4986	)	,
(	4986	)	,
(	4987	)	,
(	4988	)	,
(	4989	)	,
(	4989	)	,
(	4990	)	,
(	4991	)	,
(	4991	)	,
(	4992	)	,
(	4993	)	,
(	4994	)	,
(	4994	)	,
(	4995	)	,
(	4996	)	,
(	4996	)	,
(	4997	)	,
(	4998	)	,
(	4998	)	,
(	4999	)	,
(	5000	)	,
(	5001	)	,
(	5001	)	,
(	5002	)	,
(	5003	)	,
(	5003	)	,
(	5004	)	,
(	5005	)	,
(	5006	)	,
(	5006	)	,
(	5007	)	,
(	5008	)	,
(	5008	)	,
(	5009	)	,
(	5010	)	,
(	5010	)	,
(	5011	)	,
(	5012	)	,
(	5013	)	,
(	5013	)	,
(	5014	)	,
(	5015	)	,
(	5015	)	,
(	5016	)	,
(	5017	)	,
(	5018	)	,
(	5018	)	,
(	5019	)	,
(	5020	)	,
(	5020	)	,
(	5021	)	,
(	5022	)	,
(	5022	)	,
(	5023	)	,
(	5024	)	,
(	5025	)	,
(	5025	)	,
(	5026	)	,
(	5027	)	,
(	5027	)	,
(	5028	)	,
(	5029	)	,
(	5029	)	,
(	5030	)	,
(	5031	)	,
(	5031	)	,
(	5032	)	,
(	5033	)	,
(	5034	)	,
(	5034	)	,
(	5035	)	,
(	5036	)	,
(	5036	)	,
(	5037	)	,
(	5038	)	,
(	5038	)	,
(	5039	)	,
(	5040	)	,
(	5041	)	,
(	5041	)	,
(	5042	)	,
(	5043	)	,
(	5043	)	,
(	5044	)	,
(	5045	)	,
(	5045	)	,
(	5046	)	,
(	5047	)	,
(	5047	)	,
(	5048	)	,
(	5049	)	,
(	5050	)	,
(	5050	)	,
(	5051	)	,
(	5052	)	,
(	5052	)	,
(	5053	)	,
(	5054	)	,
(	5054	)	,
(	5055	)	,
(	5056	)	,
(	5056	)	,
(	5057	)	,
(	5058	)	,
(	5058	)	,
(	5059	)	,
(	5060	)	,
(	5061	)	,
(	5061	)	,
(	5062	)	,
(	5063	)	,
(	5063	)	,
(	5064	)	,
(	5065	)	,
(	5065	)	,
(	5066	)	,
(	5067	)	,
(	5067	)	,
(	5068	)	,
(	5069	)	,
(	5069	)	,
(	5070	)	,
(	5071	)	,
(	5071	)	,
(	5072	)	,
(	5073	)	,
(	5074	)	,
(	5074	)	,
(	5075	)	,
(	5076	)	,
(	5076	)	,
(	5077	)	,
(	5078	)	,
(	5078	)	,
(	5079	)	,
(	5080	)	,
(	5080	)	,
(	5081	)	,
(	5082	)	,
(	5082	)	,
(	5083	)	,
(	5084	)	,
(	5084	)	,
(	5085	)	,
(	5086	)	,
(	5086	)	,
(	5087	)	,
(	5088	)	,
(	5089	)	,
(	5089	)	,
(	5090	)	,
(	5091	)	,
(	5091	)	,
(	5092	)	,
(	5093	)	,
(	5093	)	,
(	5094	)	,
(	5095	)	,
(	5095	)	,
(	5096	)	,
(	5097	)	,
(	5097	)	,
(	5098	)	,
(	5099	)	,
(	5099	)	,
(	5100	)	,
(	5101	)	,
(	5101	)	,
(	5102	)	,
(	5103	)	,
(	5103	)	,
(	5104	)	,
(	5105	)	,
(	5105	)	,
(	5106	)	,
(	5107	)	,
(	5107	)	,
(	5108	)	,
(	5109	)	,
(	5109	)	,
(	5110	)	,
(	5111	)	,
(	5111	)	,
(	5112	)	,
(	5113	)	,
(	5113	)	,
(	5114	)	,
(	5115	)	,
(	5115	)	,
(	5116	)	,
(	5117	)	,
(	5117	)	,
(	5118	)	,
(	5119	)	,
(	5119	)	,
(	5120	)	,
(	5121	)	,
(	5121	)	,
(	5122	)	,
(	5123	)	,
(	5123	)	,
(	5124	)	,
(	5125	)	,
(	5125	)	,
(	5126	)	,
(	5127	)	,
(	5127	)	,
(	5128	)	,
(	5129	)	,
(	5129	)	,
(	5130	)	,
(	5131	)	,
(	5131	)	,
(	5132	)	,
(	5133	)	,
(	5133	)	,
(	5134	)	,
(	5135	)	,
(	5135	)	,
(	5136	)	,
(	5137	)	,
(	5137	)	,
(	5138	)	,
(	5139	)	,
(	5139	)	,
(	5140	)	,
(	5141	)	,
(	5141	)	,
(	5142	)	,
(	5143	)	,
(	5143	)	,
(	5144	)	,
(	5145	)	,
(	5145	)	,
(	5146	)	,
(	5147	)	,
(	5147	)	,
(	5148	)	,
(	5149	)	,
(	5149	)	,
(	5150	)	,
(	5151	)	,
(	5151	)	,
(	5152	)	,
(	5153	)	,
(	5153	)	,
(	5154	)	,
(	5155	)	,
(	5155	)	,
(	5156	)	,
(	5157	)	,
(	5157	)	,
(	5158	)	,
(	5159	)	,
(	5159	)	,
(	5160	)	,
(	5161	)	,
(	5161	)	,
(	5162	)	,
(	5162	)	,
(	5163	)	,
(	5164	)	,
(	5164	)	,
(	5165	)	,
(	5166	)	,
(	5166	)	,
(	5167	)	,
(	5168	)	,
(	5168	)	,
(	5169	)	,
(	5170	)	,
(	5170	)	,
(	5171	)	,
(	5172	)	,
(	5172	)	,
(	5173	)	,
(	5174	)	,
(	5174	)	,
(	5175	)	,
(	5176	)	,
(	5176	)	,
(	5177	)	,
(	5177	)	,
(	5178	)	,
(	5179	)	,
(	5179	)	,
(	5180	)	,
(	5181	)	,
(	5181	)	,
(	5182	)	,
(	5183	)	,
(	5183	)	,
(	5184	)	,
(	5185	)	,
(	5185	)	,
(	5186	)	,
(	5187	)	,
(	5187	)	,
(	5188	)	,
(	5188	)	,
(	5189	)	,
(	5190	)	,
(	5190	)	,
(	5191	)	,
(	5192	)	,
(	5192	)	,
(	5193	)	,
(	5194	)	,
(	5194	)	,
(	5195	)	,
(	5196	)	,
(	5196	)	,
(	5197	)	,
(	5198	)	,
(	5198	)	,
(	5199	)	,
(	5199	)	,
(	5200	)	,
(	5201	)	,
(	5201	)	,
(	5202	)	,
(	5203	)	,
(	5203	)	,
(	5204	)	,
(	5205	)	,
(	5205	)	,
(	5206	)	,
(	5207	)	,
(	5207	)	,
(	5208	)	,
(	5208	)	,
(	5209	)	,
(	5210	)	,
(	5210	)	,
(	5211	)	,
(	5212	)	,
(	5212	)	,
(	5213	)	,
(	5214	)	,
(	5214	)	,
(	5215	)	,
(	5215	)	,
(	5216	)	,
(	5217	)	,
(	5217	)	,
(	5218	)	,
(	5219	)	,
(	5219	)	,
(	5220	)	,
(	5221	)	,
(	5221	)	,
(	5222	)	,
(	5223	)	,
(	5223	)	,
(	5224	)	,
(	5224	)	,
(	5225	)	,
(	5226	)	,
(	5226	)	,
(	5227	)	,
(	5228	)	,
(	5228	)	,
(	5229	)	,
(	5229	)	,
(	5230	)	,
(	5231	)	,
(	5231	)	,
(	5232	)	,
(	5233	)	,
(	5233	)	,
(	5234	)	,
(	5235	)	,
(	5235	)	,
(	5236	)	,
(	5236	)	,
(	5237	)	,
(	5238	)	,
(	5238	)	,
(	5239	)	,
(	5240	)	,
(	5240	)	,
(	5241	)	,
(	5242	)	,
(	5242	)	,
(	5243	)	,
(	5243	)	,
(	5244	)	,
(	5245	)	,
(	5245	)	,
(	5246	)	,
(	5247	)	,
(	5247	)	,
(	5248	)	,
(	5248	)	,
(	5249	)	,
(	5250	)	,
(	5250	)	,
(	5251	)	,
(	5252	)	,
(	5252	)	,
(	5253	)	,
(	5253	)	,
(	5254	)	,
(	5255	)	,
(	5255	)	,
(	5256	)	,
(	5257	)	,
(	5257	)	,
(	5258	)	,
(	5258	)	,
(	5259	)	,
(	5260	)	,
(	5260	)	,
(	5261	)	,
(	5262	)	,
(	5262	)	,
(	5263	)	,
(	5263	)	,
(	5264	)	,
(	5265	)	,
(	5265	)	,
(	5266	)	,
(	5267	)	,
(	5267	)	,
(	5268	)	,
(	5268	)	,
(	5269	)	,
(	5270	)	,
(	5270	)	,
(	5271	)	,
(	5272	)	,
(	5272	)	,
(	5273	)	,
(	5273	)	,
(	5274	)	,
(	5275	)	,
(	5275	)	,
(	5276	)	,
(	5277	)	,
(	5277	)	,
(	5278	)	,
(	5278	)	,
(	5279	)	,
(	5280	)	,
(	5280	)	,
(	5281	)	,
(	5282	)	,
(	5282	)	,
(	5283	)	,
(	5283	)	,
(	5284	)	,
(	5285	)	,
(	5285	)	,
(	5286	)	,
(	5286	)	,
(	5287	)	,
(	5288	)	,
(	5288	)	,
(	5289	)	,
(	5290	)	,
(	5290	)	,
(	5291	)	,
(	5291	)	,
(	5292	)	,
(	5293	)	,
(	5293	)	,
(	5294	)	,
(	5294	)	,
(	5295	)	,
(	5296	)	,
(	5296	)	,
(	5297	)	,
(	5298	)	,
(	5298	)	,
(	5299	)	,
(	5299	)	,
(	5300	)	,
(	5301	)	,
(	5301	)	,
(	5302	)	,
(	5302	)	,
(	5303	)	,
(	5304	)	,
(	5304	)	,
(	5305	)	,
(	5306	)	,
(	5306	)	,
(	5307	)	,
(	5307	)	,
(	5308	)	,
(	5309	)	,
(	5309	)	,
(	5310	)	,
(	5310	)	,
(	5311	)	,
(	5312	)	,
(	5312	)	,
(	5313	)	,
(	5313	)	,
(	5314	)	,
(	5315	)	,
(	5315	)	,
(	5316	)	,
(	5317	)	,
(	5317	)	,
(	5318	)	,
(	5318	)	,
(	5319	)	,
(	5320	)	,
(	5320	)	,
(	5321	)	,
(	5321	)	,
(	5322	)	,
(	5323	)	,
(	5323	)	,
(	5324	)	,
(	5324	)	,
(	5325	)	,
(	5326	)	,
(	5326	)	,
(	5327	)	,
(	5327	)	,
(	5328	)	,
(	5329	)	,
(	5329	)	,
(	5330	)	,
(	5330	)	,
(	5331	)	,
(	5332	)	,
(	5332	)	,
(	5333	)	,
(	5333	)	,
(	5334	)	,
(	5335	)	,
(	5335	)	,
(	5336	)	,
(	5337	)	,
(	5337	)	,
(	5338	)	,
(	5338	)	,
(	5339	)	,
(	5340	)	,
(	5340	)	,
(	5341	)	,
(	5341	)	,
(	5342	)	,
(	5343	)	,
(	5343	)	,
(	5344	)	,
(	5344	)	,
(	5345	)	,
(	5346	)	,
(	5346	)	,
(	5347	)	,
(	5347	)	,
(	5348	)	,
(	5349	)	,
(	5349	)	,
(	5350	)	,
(	5350	)	,
(	5351	)	,
(	5352	)	,
(	5352	)	,
(	5353	)	,
(	5353	)	,
(	5354	)	,
(	5355	)	,
(	5355	)	,
(	5356	)	,
(	5356	)	,
(	5357	)	,
(	5358	)	,
(	5358	)	,
(	5359	)	,
(	5359	)	,
(	5360	)	,
(	5360	)	,
(	5361	)	,
(	5362	)	,
(	5362	)	,
(	5363	)	,
(	5363	)	,
(	5364	)	,
(	5365	)	,
(	5365	)	,
(	5366	)	,
(	5366	)	,
(	5367	)	,
(	5368	)	,
(	5368	)	,
(	5369	)	,
(	5369	)	,
(	5370	)	,
(	5371	)	,
(	5371	)	,
(	5372	)	,
(	5372	)	,
(	5373	)	,
(	5374	)	,
(	5374	)	,
(	5375	)	,
(	5375	)	,
(	5376	)	,
(	5377	)	,
(	5377	)	,
(	5378	)	,
(	5378	)	,
(	5379	)	,
(	5379	)	,
(	5380	)	,
(	5381	)	,
(	5381	)	,
(	5382	)	,
(	5382	)	,
(	5383	)	,
(	5384	)	,
(	5384	)	,
(	5385	)	,
(	5385	)	,
(	5386	)	,
(	5387	)	,
(	5387	)	,
(	5388	)	,
(	5388	)	,
(	5389	)	,
(	5390	)	,
(	5390	)	,
(	5391	)	,
(	5391	)	,
(	5392	)	,
(	5392	)	,
(	5393	)	,
(	5394	)	,
(	5394	)	,
(	5395	)	,
(	5395	)	,
(	5396	)	,
(	5397	)	,
(	5397	)	,
(	5398	)	,
(	5398	)	,
(	5399	)	,
(	5399	)	,
(	5400	)	,
(	5401	)	,
(	5401	)	,
(	5402	)	,
(	5402	)	,
(	5403	)	,
(	5404	)	,
(	5404	)	,
(	5405	)	,
(	5405	)	,
(	5406	)	,
(	5407	)	,
(	5407	)	,
(	5408	)	,
(	5408	)	,
(	5409	)	,
(	5409	)	,
(	5410	)	,
(	5411	)	,
(	5411	)	,
(	5412	)	,
(	5412	)	,
(	5413	)	,
(	5413	)	,
(	5414	)	,
(	5415	)	,
(	5415	)	,
(	5416	)	,
(	5416	)	,
(	5417	)	,
(	5418	)	,
(	5418	)	,
(	5419	)	,
(	5419	)	,
(	5420	)	,
(	5420	)	,
(	5421	)	,
(	5422	)	,
(	5422	)	,
(	5423	)	,
(	5423	)	,
(	5424	)	,
(	5425	)	,
(	5425	)	,
(	5426	)	,
(	5426	)	,
(	5427	)	,
(	5427	)	,
(	5428	)	,
(	5429	)	,
(	5429	)	,
(	5430	)	,
(	5430	)	,
(	5431	)	,
(	5431	)	,
(	5432	)	,
(	5433	)	,
(	5433	)	,
(	5434	)	,
(	5434	)	,
(	5435	)	,
(	5435	)	,
(	5436	)	,
(	5437	)	,
(	5437	)	,
(	5438	)	,
(	5438	)	,
(	5439	)	,
(	5440	)	,
(	5440	)	,
(	5441	)	,
(	5441	)	,
(	5442	)	,
(	5442	)	,
(	5443	)	,
(	5444	)	,
(	5444	)	,
(	5445	)	,
(	5445	)	,
(	5446	)	,
(	5446	)	,
(	5447	)	,
(	5448	)	,
(	5448	)	,
(	5449	)	,
(	5449	)	,
(	5450	)	,
(	5450	)	,
(	5451	)	,
(	5452	)	,
(	5452	)	,
(	5453	)	,
(	5453	)	,
(	5454	)	,
(	5454	)	,
(	5455	)	,
(	5456	)	,
(	5456	)	,
(	5457	)	,
(	5457	)	,
(	5458	)	,
(	5458	)	,
(	5459	)	,
(	5460	)	,
(	5460	)	,
(	5461	)	,
(	5461	)	,
(	5462	)	,
(	5462	)	,
(	5463	)	,
(	5464	)	,
(	5464	)	,
(	5465	)	,
(	5465	)	,
(	5466	)	,
(	5466	)	,
(	5467	)	,
(	5467	)	,
(	5468	)	,
(	5469	)	,
(	5469	)	,
(	5470	)	,
(	5470	)	,
(	5471	)	,
(	5471	)	,
(	5472	)	,
(	5473	)	,
(	5473	)	,
(	5474	)	,
(	5474	)	,
(	5475	)	,
(	5475	)	,
(	5476	)	,
(	5477	)	,
(	5477	)	,
(	5478	)	,
(	5478	)	,
(	5479	)	,
(	5479	)	,
(	5480	)	,
(	5480	)	,
(	5481	)	,
(	5482	)	,
(	5482	)	,
(	5483	)	,
(	5483	)	,
(	5484	)	,
(	5484	)	,
(	5485	)	,
(	5486	)	,
(	5486	)	,
(	5487	)	,
(	5487	)	,
(	5488	)	,
(	5488	)	,
(	5489	)	,
(	5489	)	,
(	5490	)	,
(	5491	)	,
(	5491	)	,
(	5492	)	,
(	5492	)	,
(	5493	)	,
(	5493	)	,
(	5494	)	,
(	5495	)	,
(	5495	)	,
(	5496	)	,
(	5496	)	,
(	5497	)	,
(	5497	)	,
(	5498	)	,
(	5498	)	,
(	5499	)	,
(	5500	)	,
(	5500	)	,
(	5501	)	,
(	5501	)	,
(	5502	)	,
(	5502	)	,
(	5503	)	,
(	5503	)	,
(	5504	)	,
(	5505	)	,
(	5505	)	,
(	5506	)	,
(	5506	)	,
(	5507	)	,
(	5507	)	,
(	5508	)	,
(	5508	)	,
(	5509	)	,
(	5510	)	,
(	5510	)	,
(	5511	)	,
(	5511	)	,
(	5512	)	,
(	5512	)	,
(	5513	)	,
(	5513	)	,
(	5514	)	,
(	5515	)	,
(	5515	)	,
(	5516	)	,
(	5516	)	,
(	5517	)	,
(	5517	)	,
(	5518	)	,
(	5518	)	,
(	5519	)	,
(	5520	)	,
(	5520	)	,
(	5521	)	,
(	5521	)	,
(	5522	)	,
(	5522	)	,
(	5523	)	,
(	5523	)	,
(	5524	)	,
(	5525	)	,
(	5525	)	,
(	5526	)	,
(	5526	)	,
(	5527	)	,
(	5527	)	,
(	5528	)	,
(	5528	)	,
(	5529	)	,
(	5530	)	,
(	5530	)	,
(	5531	)	,
(	5531	)	,
(	5532	)	,
(	5532	)	,
(	5533	)	,
(	5533	)	,
(	5534	)	,
(	5534	)	,
(	5535	)	,
(	5536	)	,
(	5536	)	,
(	5537	)	,
(	5537	)	,
(	5538	)	,
(	5538	)	,
(	5539	)	,
(	5539	)	,
(	5540	)	,
(	5540	)	,
(	5541	)	,
(	5542	)	,
(	5542	)	,
(	5543	)	,
(	5543	)	,
(	5544	)	,
(	5544	)	,
(	5545	)	,
(	5545	)	,
(	5546	)	,
(	5547	)	,
(	5547	)	,
(	5548	)	,
(	5548	)	,
(	5549	)	,
(	5549	)	,
(	5550	)	,
(	5550	)	,
(	5551	)	,
(	5551	)	,
(	5552	)	,
(	5553	)	,
(	5553	)	,
(	5554	)	,
(	5554	)	,
(	5555	)	,
(	5555	)	,
(	5556	)	,
(	5556	)	,
(	5557	)	,
(	5557	)	,
(	5558	)	,
(	5559	)	,
(	5559	)	,
(	5560	)	,
(	5560	)	,
(	5561	)	,
(	5561	)	,
(	5562	)	,
(	5562	)	,
(	5563	)	,
(	5563	)	,
(	5564	)	,
(	5564	)	,
(	5565	)	,
(	5566	)	,
(	5566	)	,
(	5567	)	,
(	5567	)	,
(	5568	)	,
(	5568	)	,
(	5569	)	,
(	5569	)	,
(	5570	)	,
(	5570	)	,
(	5571	)	,
(	5571	)	,
(	5572	)	,
(	5573	)	,
(	5573	)	,
(	5574	)	,
(	5574	)	,
(	5575	)	,
(	5575	)	,
(	5576	)	,
(	5576	)	,
(	5577	)	,
(	5577	)	,
(	5578	)	,
(	5579	)	,
(	5579	)	,
(	5580	)	,
(	5580	)	,
(	5581	)	,
(	5581	)	,
(	5582	)	,
(	5582	)	,
(	5583	)	,
(	5583	)	,
(	5584	)	,
(	5584	)	,
(	5585	)	,
(	5585	)	,
(	5586	)	,
(	5587	)	,
(	5587	)	,
(	5588	)	,
(	5588	)	,
(	5589	)	,
(	5589	)	,
(	5590	)	,
(	5590	)	,
(	5591	)	,
(	5591	)	,
(	5592	)	,
(	5592	)	,
(	5593	)	,
(	5594	)	,
(	5594	)	,
(	5595	)	,
(	5595	)	,
(	5596	)	,
(	5596	)	,
(	5597	)	,
(	5597	)	,
(	5598	)	,
(	5598	)	,
(	5599	)	,
(	5599	)	,
(	5600	)	,
(	5600	)	,
(	5601	)	,
(	5602	)	,
(	5602	)	,
(	5603	)	,
(	5603	)	,
(	5604	)	,
(	5604	)	,
(	5605	)	,
(	5605	)	,
(	5606	)	,
(	5606	)	,
(	5607	)	,
(	5607	)	,
(	5608	)	,
(	5608	)	,
(	5609	)	,
(	5609	)	,
(	5610	)	,
(	5611	)	,
(	5611	)	,
(	5612	)	,
(	5612	)	,
(	5613	)	,
(	5613	)	,
(	5614	)	,
(	5614	)	,
(	5615	)	,
(	5615	)	,
(	5616	)	,
(	5616	)	,
(	5617	)	,
(	5617	)	,
(	5618	)	,
(	5618	)	,
(	5619	)	,
(	5620	)	,
(	5620	)	,
(	5621	)	,
(	5621	)	,
(	5622	)	,
(	5622	)	,
(	5623	)	,
(	5623	)	,
(	5624	)	,
(	5624	)	,
(	5625	)	,
(	5625	)	,
(	5626	)	,
(	5626	)	,
(	5627	)	,
(	5627	)	,
(	5628	)	,
(	5628	)	,
(	5629	)	,
(	5630	)	,
(	5630	)	,
(	5631	)	,
(	5631	)	,
(	5632	)	,
(	5632	)	,
(	5633	)	,
(	5633	)	,
(	5634	)	,
(	5634	)	,
(	5635	)	,
(	5635	)	,
(	5636	)	,
(	5636	)	,
(	5637	)	,
(	5637	)	,
(	5638	)	,
(	5638	)	,
(	5639	)	,
(	5640	)	,
(	5640	)	,
(	5641	)	,
(	5641	)	,
(	5642	)	,
(	5642	)	,
(	5643	)	,
(	5643	)	,
(	5644	)	,
(	5644	)	,
(	5645	)	,
(	5645	)	,
(	5646	)	,
(	5646	)	,
(	5647	)	,
(	5647	)	,
(	5648	)	,
(	5648	)	,
(	5649	)	,
(	5649	)	,
(	5650	)	,
(	5650	)	,
(	5651	)	,
(	5651	)	,
(	5652	)	,
(	5653	)	,
(	5653	)	,
(	5654	)	,
(	5654	)	,
(	5655	)	,
(	5655	)	,
(	5656	)	,
(	5656	)	,
(	5657	)	,
(	5657	)	,
(	5658	)	,
(	5658	)	,
(	5659	)	,
(	5659	)	,
(	5660	)	
	

);

end package LUT_buzzing_pkg;