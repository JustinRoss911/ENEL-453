library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3493	)	,
(	3486	)	,
(	3479	)	,
(	3472	)	,
(	3465	)	,
(	3459	)	,
(	3452	)	,
(	3445	)	,
(	3438	)	,
(	3431	)	,
(	3425	)	,
(	3418	)	,
(	3411	)	,
(	3405	)	,
(	3398	)	,
(	3391	)	,
(	3384	)	,
(	3378	)	,
(	3371	)	,
(	3365	)	,
(	3358	)	,
(	3351	)	,
(	3345	)	,
(	3338	)	,
(	3332	)	,
(	3325	)	,
(	3319	)	,
(	3312	)	,
(	3306	)	,
(	3299	)	,
(	3293	)	,
(	3286	)	,
(	3280	)	,
(	3273	)	,
(	3267	)	,
(	3260	)	,
(	3254	)	,
(	3248	)	,
(	3241	)	,
(	3235	)	,
(	3229	)	,
(	3222	)	,
(	3216	)	,
(	3210	)	,
(	3203	)	,
(	3197	)	,
(	3191	)	,
(	3185	)	,
(	3178	)	,
(	3172	)	,
(	3166	)	,
(	3160	)	,
(	3154	)	,
(	3147	)	,
(	3141	)	,
(	3135	)	,
(	3129	)	,
(	3123	)	,
(	3117	)	,
(	3111	)	,
(	3105	)	,
(	3099	)	,
(	3093	)	,
(	3087	)	,
(	3081	)	,
(	3075	)	,
(	3069	)	,
(	3063	)	,
(	3057	)	,
(	3051	)	,
(	3045	)	,
(	3039	)	,
(	3033	)	,
(	3027	)	,
(	3021	)	,
(	3015	)	,
(	3009	)	,
(	3003	)	,
(	2998	)	,
(	2992	)	,
(	2986	)	,
(	2980	)	,
(	2974	)	,
(	2969	)	,
(	2963	)	,
(	2957	)	,
(	2951	)	,
(	2946	)	,
(	2940	)	,
(	2934	)	,
(	2929	)	,
(	2923	)	,
(	2917	)	,
(	2912	)	,
(	2906	)	,
(	2900	)	,
(	2895	)	,
(	2889	)	,
(	2883	)	,
(	2878	)	,
(	2872	)	,
(	2867	)	,
(	2861	)	,
(	2856	)	,
(	2850	)	,
(	2845	)	,
(	2839	)	,
(	2834	)	,
(	2828	)	,
(	2823	)	,
(	2817	)	,
(	2812	)	,
(	2806	)	,
(	2801	)	,
(	2796	)	,
(	2790	)	,
(	2785	)	,
(	2780	)	,
(	2774	)	,
(	2769	)	,
(	2764	)	,
(	2758	)	,
(	2753	)	,
(	2748	)	,
(	2742	)	,
(	2737	)	,
(	2732	)	,
(	2727	)	,
(	2721	)	,
(	2716	)	,
(	2711	)	,
(	2706	)	,
(	2701	)	,
(	2695	)	,
(	2690	)	,
(	2685	)	,
(	2680	)	,
(	2675	)	,
(	2670	)	,
(	2665	)	,
(	2660	)	,
(	2654	)	,
(	2649	)	,
(	2644	)	,
(	2639	)	,
(	2634	)	,
(	2629	)	,
(	2624	)	,
(	2619	)	,
(	2614	)	,
(	2609	)	,
(	2604	)	,
(	2599	)	,
(	2594	)	,
(	2589	)	,
(	2585	)	,
(	2580	)	,
(	2575	)	,
(	2570	)	,
(	2565	)	,
(	2560	)	,
(	2555	)	,
(	2550	)	,
(	2546	)	,
(	2541	)	,
(	2536	)	,
(	2531	)	,
(	2526	)	,
(	2522	)	,
(	2517	)	,
(	2512	)	,
(	2507	)	,
(	2503	)	,
(	2498	)	,
(	2493	)	,
(	2489	)	,
(	2484	)	,
(	2479	)	,
(	2474	)	,
(	2470	)	,
(	2465	)	,
(	2461	)	,
(	2456	)	,
(	2451	)	,
(	2447	)	,
(	2442	)	,
(	2438	)	,
(	2433	)	,
(	2428	)	,
(	2424	)	,
(	2419	)	,
(	2415	)	,
(	2410	)	,
(	2406	)	,
(	2401	)	,
(	2397	)	,
(	2392	)	,
(	2388	)	,
(	2383	)	,
(	2379	)	,
(	2375	)	,
(	2370	)	,
(	2366	)	,
(	2361	)	,
(	2357	)	,
(	2353	)	,
(	2348	)	,
(	2344	)	,
(	2340	)	,
(	2335	)	,
(	2331	)	,
(	2327	)	,
(	2322	)	,
(	2318	)	,
(	2314	)	,
(	2309	)	,
(	2305	)	,
(	2301	)	,
(	2297	)	,
(	2292	)	,
(	2288	)	,
(	2284	)	,
(	2280	)	,
(	2276	)	,
(	2271	)	,
(	2267	)	,
(	2263	)	,
(	2259	)	,
(	2255	)	,
(	2251	)	,
(	2246	)	,
(	2242	)	,
(	2238	)	,
(	2234	)	,
(	2230	)	,
(	2226	)	,
(	2222	)	,
(	2218	)	,
(	2214	)	,
(	2210	)	,
(	2206	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2190	)	,
(	2186	)	,
(	2182	)	,
(	2178	)	,
(	2174	)	,
(	2170	)	,
(	2166	)	,
(	2162	)	,
(	2158	)	,
(	2154	)	,
(	2150	)	,
(	2146	)	,
(	2143	)	,
(	2139	)	,
(	2135	)	,
(	2131	)	,
(	2127	)	,
(	2123	)	,
(	2120	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2101	)	,
(	2097	)	,
(	2093	)	,
(	2089	)	,
(	2086	)	,
(	2082	)	,
(	2078	)	,
(	2074	)	,
(	2071	)	,
(	2067	)	,
(	2063	)	,
(	2060	)	,
(	2056	)	,
(	2052	)	,
(	2049	)	,
(	2045	)	,
(	2042	)	,
(	2038	)	,
(	2034	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2020	)	,
(	2016	)	,
(	2013	)	,
(	2009	)	,
(	2006	)	,
(	2002	)	,
(	1999	)	,
(	1995	)	,
(	1992	)	,
(	1988	)	,
(	1985	)	,
(	1981	)	,
(	1978	)	,
(	1974	)	,
(	1971	)	,
(	1968	)	,
(	1964	)	,
(	1961	)	,
(	1957	)	,
(	1954	)	,
(	1950	)	,
(	1947	)	,
(	1944	)	,
(	1940	)	,
(	1937	)	,
(	1934	)	,
(	1930	)	,
(	1927	)	,
(	1924	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1910	)	,
(	1907	)	,
(	1904	)	,
(	1901	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1875	)	,
(	1872	)	,
(	1868	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1856	)	,
(	1853	)	,
(	1849	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1837	)	,
(	1834	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1815	)	,
(	1812	)	,
(	1809	)	,
(	1806	)	,
(	1803	)	,
(	1800	)	,
(	1797	)	,
(	1794	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1783	)	,
(	1780	)	,
(	1777	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1762	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1748	)	,
(	1745	)	,
(	1742	)	,
(	1739	)	,
(	1736	)	,
(	1733	)	,
(	1731	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1719	)	,
(	1717	)	,
(	1714	)	,
(	1711	)	,
(	1708	)	,
(	1705	)	,
(	1703	)	,
(	1700	)	,
(	1697	)	,
(	1695	)	,
(	1692	)	,
(	1689	)	,
(	1686	)	,
(	1684	)	,
(	1681	)	,
(	1678	)	,
(	1676	)	,
(	1673	)	,
(	1670	)	,
(	1668	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1649	)	,
(	1647	)	,
(	1644	)	,
(	1642	)	,
(	1639	)	,
(	1636	)	,
(	1634	)	,
(	1631	)	,
(	1629	)	,
(	1626	)	,
(	1624	)	,
(	1621	)	,
(	1619	)	,
(	1616	)	,
(	1614	)	,
(	1611	)	,
(	1609	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1596	)	,
(	1594	)	,
(	1591	)	,
(	1589	)	,
(	1586	)	,
(	1584	)	,
(	1582	)	,
(	1579	)	,
(	1577	)	,
(	1574	)	,
(	1572	)	,
(	1570	)	,
(	1567	)	,
(	1565	)	,
(	1563	)	,
(	1560	)	,
(	1558	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1548	)	,
(	1546	)	,
(	1544	)	,
(	1542	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1523	)	,
(	1521	)	,
(	1519	)	,
(	1517	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1499	)	,
(	1497	)	,
(	1495	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1412	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1405	)	,
(	1403	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1391	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1382	)	,
(	1380	)	,
(	1378	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1368	)	,
(	1366	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1344	)	,
(	1343	)	,
(	1341	)	,
(	1339	)	,
(	1338	)	,
(	1336	)	,
(	1334	)	,
(	1332	)	,
(	1331	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1322	)	,
(	1321	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1307	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1295	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1253	)	,
(	1252	)	,
(	1250	)	,
(	1249	)	,
(	1247	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	362	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	377	)	,
(	377	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	381	)	,
(	381	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	383	)	,
(	383	)	,
(	384	)	,
(	384	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	386	)	,
(	386	)	,
(	387	)	,
(	387	)	,
(	388	)	,
(	388	)	,
(	389	)	,
(	389	)	,
(	390	)	,
(	390	)	,
(	391	)	,
(	391	)	,
(	392	)	,
(	392	)	,
(	393	)	,
(	393	)	,
(	394	)	,
(	394	)	,
(	395	)	,
(	395	)	,
(	396	)	,
(	396	)	,
(	397	)	,
(	397	)	,
(	398	)	,
(	399	)	,
(	399	)	,
(	400	)	,
(	400	)	,
(	401	)	,
(	401	)	,
(	402	)	,
(	403	)	,
(	403	)	,
(	404	)	,
(	404	)	,
(	405	)	,
(	406	)	,
(	406	)	,
(	407	)	,
(	407	)	,
(	408	)	,
(	409	)	,
(	409	)	,
(	410	)	,
(	411	)	,
(	411	)	,
(	412	)	,
(	413	)	,
(	413	)	,
(	414	)	,
(	415	)	,
(	415	)	,
(	416	)	,
(	417	)	,
(	418	)	,
(	418	)	,
(	419	)	,
(	420	)	,
(	420	)	,
(	421	)	,
(	422	)	,
(	423	)	,
(	423	)	,
(	424	)	,
(	425	)	,
(	426	)	,
(	426	)	,
(	427	)	,
(	428	)	,
(	429	)	,
(	430	)	,
(	430	)	,
(	431	)	,
(	432	)	,
(	433	)	,
(	434	)	,
(	434	)	,
(	435	)	,
(	436	)	,
(	437	)	,
(	438	)	,
(	439	)	,
(	440	)	,
(	440	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	444	)	,
(	445	)	,
(	446	)	,
(	447	)	,
(	448	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	451	)	,
(	452	)	,
(	453	)	,
(	454	)	,
(	455	)	,
(	456	)	,
(	457	)	,
(	458	)	,
(	459	)	,
(	460	)	,
(	461	)	,
(	462	)	,
(	463	)	,
(	464	)	,
(	465	)	,
(	466	)	,
(	467	)	,
(	468	)	,
(	469	)	,
(	470	)	,
(	471	)	,
(	472	)	,
(	473	)	,
(	474	)	,
(	475	)	,
(	476	)	,
(	477	)	,
(	479	)	,
(	480	)	,
(	481	)	,
(	482	)	,
(	483	)	,
(	484	)	,
(	485	)	,
(	486	)	,
(	487	)	,
(	489	)	,
(	490	)	,
(	491	)	,
(	492	)	,
(	493	)	,
(	494	)	,
(	496	)	,
(	497	)	,
(	498	)	,
(	499	)	,
(	500	)	,
(	502	)	,
(	503	)	,
(	504	)	,
(	505	)	,
(	506	)	,
(	508	)	,
(	509	)	,
(	510	)	,
(	511	)	,
(	513	)	,
(	514	)	,
(	515	)	,
(	517	)	,
(	518	)	,
(	519	)	,
(	520	)	,
(	522	)	,
(	523	)	,
(	524	)	,
(	526	)	,
(	527	)	,
(	528	)	,
(	530	)	,
(	531	)	,
(	533	)	,
(	534	)	,
(	535	)	,
(	537	)	,
(	538	)	,
(	539	)	,
(	541	)	,
(	542	)	,
(	544	)	,
(	545	)	,
(	547	)	,
(	548	)	,
(	549	)	,
(	551	)	,
(	552	)	,
(	554	)	,
(	555	)	,
(	557	)	,
(	558	)	,
(	560	)	,
(	561	)	,
(	563	)	,
(	564	)	,
(	566	)	,
(	567	)	,
(	569	)	,
(	570	)	,
(	572	)	,
(	574	)	,
(	575	)	,
(	577	)	,
(	578	)	,
(	580	)	,
(	581	)	,
(	583	)	,
(	585	)	,
(	586	)	,
(	588	)	,
(	590	)	,
(	591	)	,
(	593	)	,
(	594	)	,
(	596	)	,
(	598	)	,
(	599	)	,
(	601	)	,
(	603	)	,
(	605	)	,
(	606	)	,
(	608	)	,
(	610	)	,
(	611	)	,
(	613	)	,
(	615	)	,
(	617	)	,
(	618	)	,
(	620	)	,
(	622	)	,
(	624	)	,
(	625	)	,
(	627	)	,
(	629	)	,
(	631	)	,
(	633	)	,
(	635	)	,
(	636	)	,
(	638	)	,
(	640	)	,
(	642	)	,
(	644	)	,
(	646	)	,
(	647	)	,
(	649	)	,
(	651	)	,
(	653	)	,
(	655	)	,
(	657	)	,
(	659	)	,
(	661	)	,
(	663	)	,
(	665	)	,
(	667	)	,
(	669	)	,
(	671	)	,
(	673	)	,
(	675	)	,
(	677	)	,
(	679	)	,
(	681	)	,
(	683	)	,
(	685	)	,
(	687	)	,
(	689	)	,
(	691	)	,
(	693	)	,
(	695	)	,
(	697	)	,
(	699	)	,
(	701	)	,
(	703	)	,
(	705	)	,
(	707	)	,
(	710	)	,
(	712	)	,
(	714	)	,
(	716	)	,
(	718	)	,
(	720	)	,
(	722	)	,
(	725	)	,
(	727	)	,
(	729	)	,
(	731	)	,
(	733	)	,
(	736	)	,
(	738	)	,
(	740	)	,
(	742	)	,
(	745	)	,
(	747	)	,
(	749	)	,
(	751	)	,
(	754	)	,
(	756	)	,
(	758	)	,
(	761	)	,
(	763	)	,
(	765	)	,
(	768	)	,
(	770	)	,
(	772	)	,
(	775	)	,
(	777	)	,
(	779	)	,
(	782	)	,
(	784	)	,
(	787	)	,
(	789	)	,
(	791	)	,
(	794	)	,
(	796	)	,
(	799	)	,
(	801	)	,
(	804	)	,
(	806	)	,
(	809	)	,
(	811	)	,
(	814	)	,
(	816	)	,
(	819	)	,
(	821	)	,
(	824	)	,
(	826	)	,
(	829	)	,
(	831	)	,
(	834	)	,
(	837	)	,
(	839	)	,
(	842	)	,
(	844	)	,
(	847	)	,
(	850	)	,
(	852	)	,
(	855	)	,
(	858	)	,
(	860	)	,
(	863	)	,
(	866	)	,
(	868	)	,
(	871	)	,
(	874	)	,
(	876	)	,
(	879	)	,
(	882	)	,
(	885	)	,
(	887	)	,
(	890	)	,
(	893	)	,
(	896	)	,
(	899	)	,
(	901	)	,
(	904	)	,
(	907	)	,
(	910	)	,
(	913	)	,
(	916	)	,
(	918	)	,
(	921	)	,
(	924	)	,
(	927	)	,
(	930	)	,
(	933	)	,
(	936	)	,
(	939	)	,
(	942	)	,
(	945	)	,
(	948	)	,
(	951	)	,
(	954	)	,
(	957	)	,
(	960	)	,
(	963	)	,
(	966	)	,
(	969	)	,
(	972	)	,
(	975	)	,
(	978	)	,
(	981	)	,
(	984	)	,
(	987	)	,
(	990	)	,
(	993	)	,
(	996	)	,
(	999	)	,
(	1003	)	,
(	1006	)	,
(	1009	)	,
(	1012	)	,
(	1015	)	,
(	1018	)	,
(	1022	)	,
(	1025	)	,
(	1028	)	,
(	1031	)	,
(	1035	)	,
(	1038	)	,
(	1041	)	,
(	1044	)	,
(	1048	)	,
(	1051	)	,
(	1054	)	,
(	1058	)	,
(	1061	)	,
(	1064	)	,
(	1067	)	,
(	1071	)	,
(	1074	)	,
(	1078	)	,
(	1081	)	,
(	1084	)	,
(	1088	)	,
(	1091	)	,
(	1095	)	,
(	1098	)	,
(	1101	)	,
(	1105	)	,
(	1108	)	,
(	1112	)	,
(	1115	)	,
(	1119	)	,
(	1122	)	,
(	1126	)	,
(	1129	)	,
(	1133	)	,
(	1137	)	,
(	1140	)	,
(	1144	)	,
(	1147	)	,
(	1151	)	,
(	1154	)	,
(	1158	)	,
(	1162	)	,
(	1165	)	,
(	1169	)	,
(	1173	)	,
(	1176	)	,
(	1180	)	,
(	1184	)	,
(	1187	)	,
(	1191	)	,
(	1195	)	,
(	1199	)	,
(	1202	)	,
(	1206	)	,
(	1210	)	,
(	1214	)	,
(	1217	)	,
(	1221	)	,
(	1225	)	,
(	1229	)	,
(	1233	)	,
(	1237	)	,
(	1240	)	,
(	1244	)	,
(	1248	)	,
(	1252	)	,
(	1256	)	,
(	1260	)	,
(	1264	)	,
(	1268	)	,
(	1272	)	,
(	1276	)	,
(	1280	)	,
(	1284	)	,
(	1288	)	,
(	1292	)	,
(	1296	)	,
(	1300	)	,
(	1304	)	,
(	1308	)	,
(	1312	)	,
(	1316	)	,
(	1320	)	,
(	1324	)	,
(	1328	)	,
(	1332	)	,
(	1336	)	,
(	1341	)	,
(	1345	)	,
(	1349	)	,
(	1353	)	,
(	1357	)	,
(	1362	)	,
(	1366	)	,
(	1370	)	,
(	1374	)	,
(	1378	)	,
(	1383	)	,
(	1387	)	,
(	1391	)	,
(	1396	)	,
(	1400	)	,
(	1404	)	,
(	1409	)	,
(	1413	)	,
(	1417	)	,
(	1422	)	,
(	1426	)	,
(	1430	)	,
(	1435	)	,
(	1439	)	,
(	1444	)	,
(	1448	)	,
(	1453	)	,
(	1457	)	,
(	1461	)	,
(	1466	)	,
(	1470	)	,
(	1475	)	,
(	1480	)	,
(	1484	)	,
(	1489	)	,
(	1493	)	,
(	1498	)	,
(	1502	)	,
(	1507	)	,
(	1512	)	,
(	1516	)	,
(	1521	)	,
(	1526	)	,
(	1530	)	,
(	1535	)	,
(	1540	)	,
(	1544	)	,
(	1549	)	,
(	1554	)	,
(	1558	)	,
(	1563	)	,
(	1568	)	,
(	1573	)	,
(	1578	)	,
(	1582	)	,
(	1587	)	,
(	1592	)	,
(	1597	)	,
(	1602	)	,
(	1607	)	,
(	1611	)	,
(	1616	)	,
(	1621	)	,
(	1626	)	,
(	1631	)	,
(	1636	)	,
(	1641	)	,
(	1646	)	,
(	1651	)	,
(	1656	)	,
(	1661	)	,
(	1666	)	,
(	1671	)	,
(	1676	)	,
(	1681	)	,
(	1686	)	,
(	1691	)	,
(	1696	)	,
(	1701	)	,
(	1707	)	,
(	1712	)	,
(	1717	)	,
(	1722	)	,
(	1727	)	,
(	1732	)	,
(	1738	)	,
(	1743	)	,
(	1748	)	,
(	1753	)	,
(	1759	)	,
(	1764	)	,
(	1769	)	,
(	1774	)	,
(	1780	)	,
(	1785	)	,
(	1790	)	,
(	1796	)	,
(	1801	)	,
(	1807	)	,
(	1812	)	,
(	1817	)	,
(	1823	)	,
(	1828	)	,
(	1834	)	,
(	1839	)	,
(	1845	)	,
(	1850	)	,
(	1856	)	,
(	1861	)	,
(	1867	)	,
(	1872	)	,
(	1878	)	,
(	1883	)	,
(	1889	)	,
(	1894	)	,
(	1900	)	,
(	1906	)	,
(	1911	)	,
(	1917	)	,
(	1923	)	,
(	1928	)	,
(	1934	)	,
(	1940	)	,
(	1946	)	,
(	1951	)	,
(	1957	)	,
(	1963	)	,
(	1969	)	,
(	1974	)	,
(	1980	)	,
(	1986	)	,
(	1992	)	,
(	1998	)	,
(	2004	)	,
(	2009	)	,
(	2015	)	,
(	2021	)	,
(	2027	)	,
(	2033	)	,
(	2039	)	,
(	2045	)	,
(	2051	)	,
(	2057	)	,
(	2063	)	,
(	2069	)	,
(	2075	)	,
(	2081	)	,
(	2087	)	,
(	2093	)	,
(	2099	)	,
(	2106	)	,
(	2112	)	,
(	2118	)	,
(	2124	)	,
(	2130	)	,
(	2136	)	,
(	2143	)	,
(	2149	)	,
(	2155	)	,
(	2161	)	,
(	2167	)	,
(	2174	)	,
(	2180	)	,
(	2186	)	,
(	2193	)	,
(	2199	)	,
(	2205	)	,
(	2212	)	,
(	2218	)	,
(	2225	)	,
(	2231	)	,
(	2237	)	,
(	2244	)	,
(	2250	)	,
(	2257	)	,
(	2263	)	,
(	2270	)	,
(	2276	)	,
(	2283	)	,
(	2289	)	,
(	2296	)	,
(	2302	)	,
(	2309	)	,
(	2316	)	,
(	2322	)	,
(	2329	)	,
(	2336	)	,
(	2342	)	,
(	2349	)	,
(	2356	)	,
(	2362	)	,
(	2369	)	,
(	2376	)	,
(	2383	)	,
(	2389	)	,
(	2396	)	,
(	2403	)	,
(	2410	)	,
(	2417	)	,
(	2423	)	,
(	2430	)	,
(	2437	)	,
(	2444	)	,
(	2451	)	,
(	2458	)	,
(	2465	)	,
(	2472	)	,
(	2479	)	,
(	2486	)	,
(	2493	)	,
(	2500	)	,
(	2507	)	,
(	2514	)	,
(	2521	)	,
(	2528	)	,
(	2535	)	,
(	2542	)	,
(	2550	)	,
(	2557	)	,
(	2564	)	,
(	2571	)	,
(	2578	)	,
(	2585	)	,
(	2593	)	,
(	2600	)	,
(	2607	)	,
(	2615	)	,
(	2622	)	,
(	2629	)	,
(	2636	)	,
(	2644	)	,
(	2651	)	,
(	2659	)	,
(	2666	)	,
(	2673	)	,
(	2681	)	,
(	2688	)	,
(	2696	)	,
(	2703	)	,
(	2711	)	,
(	2718	)	,
(	2726	)	,
(	2733	)	,
(	2741	)	,
(	2748	)	,
(	2756	)	,
(	2764	)	,
(	2771	)	,
(	2779	)	,
(	2787	)	,
(	2794	)	,
(	2802	)	,
(	2810	)	,
(	2817	)	,
(	2825	)	,
(	2833	)	,
(	2841	)	,
(	2849	)	,
(	2856	)	,
(	2864	)	,
(	2872	)	,
(	2880	)	,
(	2888	)	,
(	2896	)	,
(	2904	)	,
(	2912	)	,
(	2920	)	,
(	2927	)	,
(	2935	)	,
(	2943	)	,
(	2952	)	,
(	2960	)	,
(	2968	)	,
(	2976	)	,
(	2984	)	,
(	2992	)	,
(	3000	)	,
(	3008	)	,
(	3016	)	,
(	3024	)	,
(	3033	)	,
(	3041	)	,
(	3049	)	,
(	3057	)	,
(	3066	)	,
(	3074	)	,
(	3082	)	,
(	3091	)	,
(	3099	)	,
(	3107	)	,
(	3116	)	,
(	3124	)	,
(	3132	)	,
(	3141	)	,
(	3149	)	,
(	3158	)	,
(	3166	)	,
(	3175	)	,
(	3183	)	,
(	3192	)	,
(	3200	)	,
(	3209	)	,
(	3217	)	,
(	3226	)	,
(	3235	)	,
(	3243	)	,
(	3252	)	,
(	3261	)	,
(	3269	)	,
(	3278	)	,
(	3287	)	,
(	3295	)	,
(	3304	)	,
(	3313	)	,
(	3322	)	,
(	3331	)	,
(	3339	)	,
(	3348	)	,
(	3357	)	,
(	3366	)	,
(	3375	)	,
(	3384	)	,
(	3393	)	,
(	3402	)	,
(	3411	)	,
(	3420	)	,
(	3429	)	,
(	3438	)	,
(	3447	)	,
(	3456	)	,
(	3465	)	,
(	3474	)	,
(	3483	)	,
(	3492	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	,
(	3500	)	

);


end package LUT_pkg;
