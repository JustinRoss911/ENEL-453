library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	5414	)	, -- array index 0 (voltage = "000000000000" or 0 mV), distance output 54.14 (54.14 cm)
(	5405	)	, -- array index 1 (voltage = "000000000001" or 1 mV), distance output 54.05 (54.05 cm)
(	5396	)	,
(	5387	)	,
(	5379	)	,
(	5370	)	, -- array index 5 (voltage = "000000000101" or 5 mV), distance output 53.70 (53.70 cm)
(	5361	)	,
(	5353	)	,
(	5344	)	,
(	5336	)	,
(	5327	)	,
(	5318	)	,
(	5310	)	,
(	5301	)	,
(	5293	)	,
(	5284	)	,
(	5276	)	,
(	5267	)	,
(	5259	)	,
(	5250	)	,
(	5242	)	,
(	5233	)	,
(	5225	)	,
(	5217	)	,
(	5208	)	,
(	5200	)	,
(	5191	)	,
(	5183	)	,
(	5175	)	,
(	5166	)	,
(	5158	)	,
(	5150	)	,
(	5141	)	,
(	5133	)	,
(	5125	)	,
(	5116	)	,
(	5108	)	,
(	5100	)	,
(	5092	)	,
(	5083	)	,
(	5075	)	,
(	5067	)	,
(	5059	)	,
(	5051	)	,
(	5042	)	,
(	5034	)	,
(	5026	)	,
(	5018	)	,
(	5010	)	,
(	5002	)	,
(	4994	)	,
(	4986	)	,
(	4977	)	,
(	4969	)	,
(	4961	)	,
(	4953	)	,
(	4945	)	,
(	4937	)	,
(	4929	)	,
(	4921	)	,
(	4913	)	,
(	4905	)	,
(	4897	)	,
(	4889	)	,
(	4882	)	,
(	4874	)	,
(	4866	)	,
(	4858	)	,
(	4850	)	,
(	4842	)	,
(	4834	)	,
(	4826	)	,
(	4819	)	,
(	4811	)	,
(	4803	)	,
(	4795	)	,
(	4787	)	,
(	4780	)	,
(	4772	)	,
(	4764	)	,
(	4756	)	,
(	4749	)	,
(	4741	)	,
(	4733	)	,
(	4726	)	,
(	4718	)	,
(	4710	)	,
(	4702	)	,
(	4695	)	,
(	4687	)	,
(	4680	)	,
(	4672	)	,
(	4664	)	,
(	4657	)	,
(	4649	)	,
(	4642	)	,
(	4634	)	,
(	4627	)	,
(	4619	)	,
(	4612	)	,
(	4604	)	,
(	4597	)	,
(	4589	)	,
(	4582	)	,
(	4574	)	,
(	4567	)	,
(	4559	)	,
(	4552	)	,
(	4544	)	,
(	4537	)	,
(	4530	)	,
(	4522	)	,
(	4515	)	,
(	4507	)	,
(	4500	)	,
(	4493	)	,
(	4485	)	,
(	4478	)	,
(	4471	)	,
(	4464	)	,
(	4456	)	,
(	4449	)	,
(	4442	)	,
(	4435	)	,
(	4427	)	,
(	4420	)	,
(	4413	)	,
(	4406	)	,
(	4398	)	,
(	4391	)	,
(	4384	)	,
(	4377	)	,
(	4370	)	,
(	4363	)	,
(	4356	)	,
(	4348	)	,
(	4341	)	,
(	4334	)	,
(	4327	)	,
(	4320	)	,
(	4313	)	,
(	4306	)	,
(	4299	)	,
(	4292	)	,
(	4285	)	,
(	4278	)	,
(	4271	)	,
(	4264	)	,
(	4257	)	,
(	4250	)	,
(	4243	)	,
(	4236	)	,
(	4229	)	,
(	4222	)	,
(	4215	)	,
(	4208	)	,
(	4202	)	,
(	4195	)	,
(	4188	)	,
(	4181	)	,
(	4174	)	,
(	4167	)	,
(	4161	)	,
(	4154	)	,
(	4147	)	,
(	4140	)	,
(	4133	)	,
(	4127	)	,
(	4120	)	,
(	4113	)	,
(	4106	)	,
(	4100	)	,
(	4093	)	,
(	4086	)	,
(	4080	)	,
(	4073	)	,
(	4066	)	,
(	4060	)	,
(	4053	)	,
(	4046	)	,
(	4040	)	,
(	4033	)	,
(	4026	)	,
(	4020	)	,
(	4013	)	,
(	4007	)	,
(	4000	)	,
(	3993	)	,
(	3987	)	,
(	3980	)	,
(	3974	)	,
(	3967	)	,
(	3961	)	,
(	3954	)	,
(	3948	)	,
(	3941	)	,
(	3935	)	,
(	3929	)	,
(	3922	)	,
(	3916	)	,
(	3909	)	,
(	3903	)	,
(	3896	)	,
(	3890	)	,
(	3884	)	,
(	3877	)	,
(	3871	)	,
(	3865	)	,
(	3858	)	,
(	3852	)	,
(	3846	)	,
(	3839	)	,
(	3833	)	,
(	3827	)	,
(	3820	)	,
(	3814	)	,
(	3808	)	,
(	3802	)	,
(	3795	)	,
(	3789	)	,
(	3783	)	,
(	3777	)	,
(	3771	)	,
(	3764	)	,
(	3758	)	,
(	3752	)	,
(	3746	)	,
(	3740	)	,
(	3734	)	,
(	3727	)	,
(	3721	)	,
(	3715	)	,
(	3709	)	,
(	3703	)	,
(	3697	)	,
(	3691	)	,
(	3685	)	,
(	3679	)	,
(	3673	)	,
(	3667	)	,
(	3661	)	,
(	3655	)	,
(	3649	)	,
(	3643	)	,
(	3637	)	,
(	3631	)	,
(	3625	)	,
(	3619	)	,
(	3613	)	,
(	3607	)	,
(	3601	)	,
(	3595	)	,
(	3589	)	,
(	3583	)	,
(	3577	)	,
(	3572	)	,
(	3566	)	,
(	3560	)	,
(	3554	)	,
(	3548	)	,
(	3542	)	,
(	3537	)	,
(	3531	)	,
(	3525	)	,
(	3519	)	,
(	3513	)	,
(	3508	)	,
(	3502	)	,
(	3496	)	,
(	3490	)	,
(	3485	)	,
(	3479	)	,
(	3473	)	,
(	3468	)	,
(	3462	)	,
(	3456	)	,
(	3450	)	,
(	3445	)	,
(	3439	)	,
(	3434	)	,
(	3428	)	,
(	3422	)	,
(	3417	)	,
(	3411	)	,
(	3405	)	,
(	3400	)	,
(	3394	)	,
(	3389	)	,
(	3383	)	,
(	3378	)	,
(	3372	)	,
(	3366	)	,
(	3361	)	,
(	3355	)	,
(	3350	)	,
(	3344	)	,
(	3339	)	,
(	3333	)	,
(	3328	)	,
(	3323	)	,
(	3317	)	,
(	3312	)	,
(	3306	)	,
(	3301	)	,
(	3295	)	,
(	3290	)	,
(	3285	)	,
(	3279	)	,
(	3274	)	,
(	3268	)	,
(	3263	)	,
(	3258	)	,
(	3252	)	,
(	3247	)	,
(	3242	)	,
(	3236	)	,
(	3231	)	,
(	3226	)	,
(	3221	)	,
(	3215	)	,
(	3210	)	,
(	3205	)	,
(	3199	)	,
(	3194	)	,
(	3189	)	,
(	3184	)	,
(	3179	)	,
(	3173	)	,
(	3168	)	,
(	3163	)	,
(	3158	)	,
(	3153	)	,
(	3147	)	,
(	3142	)	,
(	3137	)	,
(	3132	)	,
(	3127	)	,
(	3122	)	,
(	3117	)	,
(	3112	)	,
(	3106	)	,
(	3101	)	,
(	3096	)	,
(	3091	)	,
(	3086	)	,
(	3081	)	,
(	3076	)	,
(	3071	)	,
(	3066	)	,
(	3061	)	,
(	3056	)	,
(	3051	)	,
(	3046	)	,
(	3041	)	,
(	3036	)	,
(	3031	)	,
(	3026	)	,
(	3021	)	,
(	3016	)	,
(	3011	)	,
(	3006	)	,
(	3001	)	,
(	2997	)	,
(	2992	)	,
(	2987	)	,
(	2982	)	,
(	2977	)	,
(	2972	)	,
(	2967	)	,
(	2962	)	,
(	2958	)	,
(	2953	)	,
(	2948	)	,
(	2943	)	,
(	2938	)	,
(	2934	)	,
(	2929	)	,
(	2924	)	,
(	2919	)	,
(	2914	)	,
(	2910	)	,
(	2905	)	,
(	2900	)	,
(	2896	)	,
(	2891	)	,
(	2886	)	,
(	2881	)	,
(	2877	)	,
(	2872	)	,
(	2867	)	,
(	2863	)	,
(	2858	)	,
(	2853	)	,
(	2849	)	,
(	2844	)	,
(	2839	)	,
(	2835	)	,
(	2830	)	,
(	2826	)	,
(	2821	)	,
(	2816	)	,
(	2812	)	,
(	2807	)	,
(	2803	)	,
(	2798	)	,
(	2794	)	,
(	2789	)	,
(	2784	)	,
(	2780	)	,
(	2775	)	,
(	2771	)	,
(	2766	)	,
(	2762	)	,
(	2757	)	,
(	2753	)	,
(	2748	)	,
(	2744	)	,
(	2740	)	,
(	2735	)	,
(	2731	)	,
(	2726	)	,
(	2722	)	,
(	2717	)	,
(	2713	)	,
(	2709	)	,
(	2704	)	,
(	2700	)	,
(	2695	)	,
(	2691	)	,
(	2687	)	,
(	2682	)	,
(	2678	)	,
(	2674	)	,
(	2669	)	,
(	2665	)	,
(	2661	)	,
(	2656	)	,
(	2652	)	,
(	2648	)	,
(	2643	)	,
(	2639	)	,
(	2635	)	,
(	2631	)	,
(	2626	)	,
(	2622	)	,
(	2618	)	,
(	2614	)	,
(	2610	)	,
(	2605	)	,
(	2601	)	,
(	2597	)	,
(	2593	)	,
(	2589	)	,
(	2584	)	,
(	2580	)	,
(	2576	)	,
(	2572	)	,
(	2568	)	,
(	2564	)	,
(	2559	)	,
(	2555	)	,
(	2551	)	,
(	2547	)	,
(	2543	)	,
(	2539	)	,
(	2535	)	,
(	2531	)	,
(	2527	)	,
(	2523	)	,
(	2518	)	,
(	2514	)	,
(	2510	)	,
(	2506	)	,
(	2502	)	,
(	2498	)	,
(	2494	)	,
(	2490	)	,
(	2486	)	,
(	2482	)	,
(	2478	)	,
(	2474	)	,
(	2470	)	,
(	2466	)	,
(	2462	)	,
(	2459	)	,
(	2455	)	,
(	2451	)	,
(	2447	)	,
(	2443	)	,
(	2439	)	,
(	2435	)	,
(	2431	)	,
(	2427	)	,
(	2423	)	,
(	2419	)	,
(	2416	)	,
(	2412	)	,
(	2408	)	,
(	2404	)	,
(	2400	)	,
(	2396	)	,
(	2392	)	,
(	2389	)	,
(	2385	)	,
(	2381	)	,
(	2377	)	,
(	2373	)	,
(	2370	)	,
(	2366	)	,
(	2362	)	,
(	2358	)	,
(	2355	)	,
(	2351	)	,
(	2347	)	,
(	2343	)	,
(	2340	)	,
(	2336	)	,
(	2332	)	,
(	2328	)	,
(	2325	)	,
(	2321	)	,
(	2317	)	,
(	2314	)	,
(	2310	)	,
(	2306	)	,
(	2303	)	,
(	2299	)	,
(	2295	)	,
(	2292	)	,
(	2288	)	,
(	2285	)	,
(	2281	)	,
(	2277	)	,
(	2274	)	,
(	2270	)	,
(	2266	)	,
(	2263	)	,
(	2259	)	,
(	2256	)	,
(	2252	)	,
(	2249	)	,
(	2245	)	,
(	2242	)	,
(	2238	)	,
(	2234	)	,
(	2231	)	,
(	2227	)	,
(	2224	)	,
(	2220	)	,
(	2217	)	,
(	2213	)	,
(	2210	)	,
(	2206	)	,
(	2203	)	,
(	2199	)	,
(	2196	)	,
(	2193	)	,
(	2189	)	,
(	2186	)	,
(	2182	)	,
(	2179	)	,
(	2175	)	,
(	2172	)	,
(	2169	)	,
(	2165	)	,
(	2162	)	,
(	2158	)	,
(	2155	)	,
(	2152	)	,
(	2148	)	,
(	2145	)	,
(	2142	)	,
(	2138	)	,
(	2135	)	,
(	2131	)	,
(	2128	)	,
(	2125	)	,
(	2122	)	,
(	2118	)	,
(	2115	)	,
(	2112	)	,
(	2108	)	,
(	2105	)	,
(	2102	)	,
(	2098	)	,
(	2095	)	,
(	2092	)	,
(	2089	)	,
(	2085	)	,
(	2082	)	,
(	2079	)	,
(	2076	)	,
(	2073	)	,
(	2069	)	,
(	2066	)	,
(	2063	)	,
(	2060	)	,
(	2056	)	,
(	2053	)	,
(	2050	)	,
(	2047	)	,
(	2044	)	,
(	2041	)	,
(	2037	)	,
(	2034	)	,
(	2031	)	,
(	2028	)	,
(	2025	)	,
(	2022	)	,
(	2019	)	,
(	2016	)	,
(	2012	)	,
(	2009	)	,
(	2006	)	,
(	2003	)	,
(	2000	)	,
(	1997	)	,
(	1994	)	,
(	1991	)	,
(	1988	)	,
(	1985	)	,
(	1982	)	,
(	1979	)	,
(	1976	)	,
(	1973	)	,
(	1970	)	,
(	1967	)	,
(	1964	)	,
(	1960	)	,
(	1957	)	,
(	1955	)	,
(	1952	)	,
(	1949	)	,
(	1946	)	,
(	1943	)	,
(	1940	)	,
(	1937	)	,
(	1934	)	,
(	1931	)	,
(	1928	)	,
(	1925	)	,
(	1922	)	,
(	1919	)	,
(	1916	)	,
(	1913	)	,
(	1910	)	,
(	1907	)	,
(	1904	)	,
(	1902	)	,
(	1899	)	,
(	1896	)	,
(	1893	)	,
(	1890	)	,
(	1887	)	,
(	1884	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1856	)	,
(	1853	)	,
(	1851	)	,
(	1848	)	,
(	1845	)	,
(	1842	)	,
(	1839	)	,
(	1837	)	,
(	1834	)	,
(	1831	)	,
(	1828	)	,
(	1826	)	,
(	1823	)	,
(	1820	)	,
(	1817	)	,
(	1815	)	,
(	1812	)	,
(	1809	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1799	)	,
(	1796	)	,
(	1793	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1783	)	,
(	1780	)	,
(	1777	)	,
(	1775	)	,
(	1772	)	,
(	1769	)	,
(	1767	)	,
(	1764	)	,
(	1762	)	,
(	1759	)	,
(	1756	)	,
(	1754	)	,
(	1751	)	,
(	1749	)	,
(	1746	)	,
(	1743	)	,
(	1741	)	,
(	1738	)	,
(	1736	)	,
(	1733	)	,
(	1731	)	,
(	1728	)	,
(	1726	)	,
(	1723	)	,
(	1721	)	,
(	1718	)	,
(	1715	)	,
(	1713	)	,
(	1710	)	,
(	1708	)	,
(	1705	)	,
(	1703	)	,
(	1700	)	,
(	1698	)	,
(	1696	)	,
(	1693	)	,
(	1691	)	,
(	1688	)	,
(	1686	)	,
(	1683	)	,
(	1681	)	,
(	1678	)	,
(	1676	)	,
(	1673	)	,
(	1671	)	,
(	1669	)	,
(	1666	)	,
(	1664	)	,
(	1661	)	,
(	1659	)	,
(	1657	)	,
(	1654	)	,
(	1652	)	,
(	1649	)	,
(	1647	)	,
(	1645	)	,
(	1642	)	,
(	1640	)	,
(	1638	)	,
(	1635	)	,
(	1633	)	,
(	1631	)	,
(	1628	)	,
(	1626	)	,
(	1624	)	,
(	1621	)	,
(	1619	)	,
(	1617	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1607	)	,
(	1605	)	,
(	1603	)	,
(	1601	)	,
(	1598	)	,
(	1596	)	,
(	1594	)	,
(	1591	)	,
(	1589	)	,
(	1587	)	,
(	1585	)	,
(	1582	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1565	)	,
(	1563	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1536	)	,
(	1534	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1519	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1499	)	,
(	1497	)	,
(	1495	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1445	)	,
(	1443	)	,
(	1441	)	,
(	1439	)	,
(	1437	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1405	)	,
(	1403	)	,
(	1401	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1382	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1373	)	,
(	1372	)	,
(	1370	)	,
(	1368	)	,
(	1366	)	,
(	1365	)	,
(	1363	)	,
(	1361	)	,
(	1359	)	,
(	1357	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1350	)	,
(	1349	)	,
(	1347	)	,
(	1345	)	,
(	1344	)	,
(	1342	)	,
(	1340	)	,
(	1338	)	,
(	1337	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1330	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1321	)	,
(	1320	)	,
(	1318	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1306	)	,
(	1305	)	,
(	1303	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1293	)	,
(	1292	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1266	)	,
(	1265	)	,
(	1263	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1234	)	,
(	1233	)	,
(	1231	)	,
(	1230	)	,
(	1228	)	,
(	1227	)	,
(	1225	)	,
(	1224	)	,
(	1223	)	,
(	1221	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1215	)	,
(	1214	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1205	)	,
(	1204	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	488	)	,
(	488	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	491	)	,
(	491	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	493	)	,
(	493	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	495	)	,
(	495	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	497	)	,
(	497	)	,
(	498	)	,
(	498	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	500	)	,
(	500	)	,
(	501	)	,
(	501	)	,
(	502	)	,
(	502	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	504	)	,
(	504	)	,
(	505	)	,
(	505	)	,
(	506	)	,
(	506	)	,
(	507	)	,
(	507	)	,
(	508	)	,
(	508	)	,
(	509	)	,
(	509	)	,
(	510	)	,
(	510	)	,
(	511	)	,
(	511	)	,
(	512	)	,
(	512	)	,
(	513	)	,
(	513	)	,
(	514	)	,
(	514	)	,
(	515	)	,
(	515	)	,
(	516	)	,
(	516	)	,
(	517	)	,
(	517	)	,
(	518	)	,
(	518	)	,
(	519	)	,
(	519	)	,
(	520	)	,
(	521	)	,
(	521	)	,
(	522	)	,
(	522	)	,
(	523	)	,
(	523	)	,
(	524	)	,
(	524	)	,
(	525	)	,
(	526	)	,
(	526	)	,
(	527	)	,
(	527	)	,
(	528	)	,
(	529	)	,
(	529	)	,
(	530	)	,
(	530	)	,
(	531	)	,
(	532	)	,
(	532	)	,
(	533	)	,
(	533	)	,
(	534	)	,
(	535	)	,
(	535	)	,
(	536	)	,
(	536	)	,
(	537	)	,
(	538	)	,
(	538	)	,
(	539	)	,
(	540	)	,
(	540	)	,
(	541	)	,
(	542	)	,
(	542	)	,
(	543	)	,
(	544	)	,
(	544	)	,
(	545	)	,
(	546	)	,
(	546	)	,
(	547	)	,
(	548	)	,
(	548	)	,
(	549	)	,
(	550	)	,
(	550	)	,
(	551	)	,
(	552	)	,
(	552	)	,
(	553	)	,
(	554	)	,
(	554	)	,
(	555	)	,
(	556	)	,
(	557	)	,
(	557	)	,
(	558	)	,
(	559	)	,
(	560	)	,
(	560	)	,
(	561	)	,
(	562	)	,
(	562	)	,
(	563	)	,
(	564	)	,
(	565	)	,
(	565	)	,
(	566	)	,
(	567	)	,
(	568	)	,
(	568	)	,
(	569	)	,
(	570	)	,
(	571	)	,
(	572	)	,
(	572	)	,
(	573	)	,
(	574	)	,
(	575	)	,
(	576	)	,
(	576	)	,
(	577	)	,
(	578	)	,
(	579	)	,
(	580	)	,
(	580	)	,
(	581	)	,
(	582	)	,
(	583	)	,
(	584	)	,
(	585	)	,
(	585	)	,
(	586	)	,
(	587	)	,
(	588	)	,
(	589	)	,
(	590	)	,
(	590	)	,
(	591	)	,
(	592	)	,
(	593	)	,
(	594	)	,
(	595	)	,
(	596	)	,
(	597	)	,
(	597	)	,
(	598	)	,
(	599	)	,
(	600	)	,
(	601	)	,
(	602	)	,
(	603	)	,
(	604	)	,
(	605	)	,
(	605	)	,
(	606	)	,
(	607	)	,
(	608	)	,
(	609	)	,
(	610	)	,
(	611	)	,
(	612	)	,
(	613	)	,
(	614	)	,
(	615	)	,
(	616	)	,
(	617	)	,
(	618	)	,
(	619	)	,
(	620	)	,
(	621	)	,
(	622	)	,
(	623	)	,
(	624	)	,
(	625	)	,
(	626	)	,
(	627	)	,
(	628	)	,
(	629	)	,
(	630	)	,
(	631	)	,
(	632	)	,
(	633	)	,
(	634	)	,
(	635	)	,
(	636	)	,
(	637	)	,
(	638	)	,
(	639	)	,
(	640	)	,
(	641	)	,
(	642	)	,
(	643	)	,
(	644	)	,
(	645	)	,
(	646	)	,
(	647	)	,
(	648	)	,
(	649	)	,
(	650	)	,
(	651	)	,
(	653	)	,
(	654	)	,
(	655	)	,
(	656	)	,
(	657	)	,
(	658	)	,
(	659	)	,
(	660	)	,
(	661	)	,
(	662	)	,
(	664	)	,
(	665	)	,
(	666	)	,
(	667	)	,
(	668	)	,
(	669	)	,
(	670	)	,
(	672	)	,
(	673	)	,
(	674	)	,
(	675	)	,
(	676	)	,
(	677	)	,
(	679	)	,
(	680	)	,
(	681	)	,
(	682	)	,
(	683	)	,
(	685	)	,
(	686	)	,
(	687	)	,
(	688	)	,
(	689	)	,
(	691	)	,
(	692	)	,
(	693	)	,
(	694	)	,
(	695	)	,
(	697	)	,
(	698	)	,
(	699	)	,
(	700	)	,
(	702	)	,
(	703	)	,
(	704	)	,
(	705	)	,
(	707	)	,
(	708	)	,
(	709	)	,
(	711	)	,
(	712	)	,
(	713	)	,
(	714	)	,
(	716	)	,
(	717	)	,
(	718	)	,
(	720	)	,
(	721	)	,
(	722	)	,
(	724	)	,
(	725	)	,
(	726	)	,
(	728	)	,
(	729	)	,
(	730	)	,
(	732	)	,
(	733	)	,
(	734	)	,
(	736	)	,
(	737	)	,
(	739	)	,
(	740	)	,
(	741	)	,
(	743	)	,
(	744	)	,
(	745	)	,
(	747	)	,
(	748	)	,
(	750	)	,
(	751	)	,
(	752	)	,
(	754	)	,
(	755	)	,
(	757	)	,
(	758	)	,
(	760	)	,
(	761	)	,
(	762	)	,
(	764	)	,
(	765	)	,
(	767	)	,
(	768	)	,
(	770	)	,
(	771	)	,
(	773	)	,
(	774	)	,
(	776	)	,
(	777	)	,
(	779	)	,
(	780	)	,
(	782	)	,
(	783	)	,
(	785	)	,
(	786	)	,
(	788	)	,
(	789	)	,
(	791	)	,
(	792	)	,
(	794	)	,
(	795	)	,
(	797	)	,
(	799	)	,
(	800	)	,
(	802	)	,
(	803	)	,
(	805	)	,
(	806	)	,
(	808	)	,
(	810	)	,
(	811	)	,
(	813	)	,
(	814	)	,
(	816	)	,
(	818	)	,
(	819	)	,
(	821	)	,
(	822	)	,
(	824	)	,
(	826	)	,
(	827	)	,
(	829	)	,
(	831	)	,
(	832	)	,
(	834	)	,
(	836	)	,
(	837	)	,
(	839	)	,
(	841	)	,
(	842	)	,
(	844	)	,
(	846	)	,
(	847	)	,
(	849	)	,
(	851	)	,
(	853	)	,
(	854	)	,
(	856	)	,
(	858	)	,
(	859	)	,
(	861	)	,
(	863	)	,
(	865	)	,
(	866	)	,
(	868	)	,
(	870	)	,
(	872	)	,
(	874	)	,
(	875	)	,
(	877	)	,
(	879	)	,
(	881	)	,
(	882	)	,
(	884	)	,
(	886	)	,
(	888	)	,
(	890	)	,
(	892	)	,
(	893	)	,
(	895	)	,
(	897	)	,
(	899	)	,
(	901	)	,
(	903	)	,
(	904	)	,
(	906	)	,
(	908	)	,
(	910	)	,
(	912	)	,
(	914	)	,
(	916	)	,
(	918	)	,
(	920	)	,
(	921	)	,
(	923	)	,
(	925	)	,
(	927	)	,
(	929	)	,
(	931	)	,
(	933	)	,
(	935	)	,
(	937	)	,
(	939	)	,
(	941	)	,
(	943	)	,
(	945	)	,
(	947	)	,
(	949	)	,
(	951	)	,
(	953	)	,
(	955	)	,
(	957	)	,
(	959	)	,
(	961	)	,
(	963	)	,
(	965	)	,
(	967	)	,
(	969	)	,
(	971	)	,
(	973	)	,
(	975	)	,
(	977	)	,
(	979	)	,
(	981	)	,
(	983	)	,
(	985	)	,
(	987	)	,
(	989	)	,
(	992	)	,
(	994	)	,
(	996	)	,
(	998	)	,
(	1000	)	,
(	1002	)	,
(	1004	)	,
(	1006	)	,
(	1008	)	,
(	1011	)	,
(	1013	)	,
(	1015	)	,
(	1017	)	,
(	1019	)	,
(	1021	)	,
(	1024	)	,
(	1026	)	,
(	1028	)	,
(	1030	)	,
(	1032	)	,
(	1035	)	,
(	1037	)	,
(	1039	)	,
(	1041	)	,
(	1043	)	,
(	1046	)	,
(	1048	)	,
(	1050	)	,
(	1052	)	,
(	1055	)	,
(	1057	)	,
(	1059	)	,
(	1061	)	,
(	1064	)	,
(	1066	)	,
(	1068	)	,
(	1071	)	,
(	1073	)	,
(	1075	)	,
(	1078	)	,
(	1080	)	,
(	1082	)	,
(	1085	)	,
(	1087	)	,
(	1089	)	,
(	1092	)	,
(	1094	)	,
(	1096	)	,
(	1099	)	,
(	1101	)	,
(	1103	)	,
(	1106	)	,
(	1108	)	,
(	1111	)	,
(	1113	)	,
(	1115	)	,
(	1118	)	,
(	1120	)	,
(	1123	)	,
(	1125	)	,
(	1128	)	,
(	1130	)	,
(	1132	)	,
(	1135	)	,
(	1137	)	,
(	1140	)	,
(	1142	)	,
(	1145	)	,
(	1147	)	,
(	1150	)	,
(	1152	)	,
(	1155	)	,
(	1157	)	,
(	1160	)	,
(	1162	)	,
(	1165	)	,
(	1167	)	,
(	1170	)	,
(	1173	)	,
(	1175	)	,
(	1178	)	,
(	1180	)	,
(	1183	)	,
(	1185	)	,
(	1188	)	,
(	1191	)	,
(	1193	)	,
(	1196	)	,
(	1198	)	,
(	1201	)	,
(	1204	)	,
(	1206	)	,
(	1209	)	,
(	1212	)	,
(	1214	)	,
(	1217	)	,
(	1220	)	,
(	1222	)	,
(	1225	)	,
(	1228	)	,
(	1230	)	,
(	1233	)	,
(	1236	)	,
(	1238	)	,
(	1241	)	,
(	1244	)	,
(	1247	)	,
(	1249	)	,
(	1252	)	,
(	1255	)	,
(	1258	)	,
(	1260	)	,
(	1263	)	,
(	1266	)	,
(	1269	)	,
(	1271	)	,
(	1274	)	,
(	1277	)	,
(	1280	)	,
(	1283	)	,
(	1285	)	,
(	1288	)	,
(	1291	)	,
(	1294	)	,
(	1297	)	,
(	1300	)	,
(	1302	)	,
(	1305	)	,
(	1308	)	,
(	1311	)	,
(	1314	)	,
(	1317	)	,
(	1320	)	,
(	1323	)	,
(	1326	)	,
(	1329	)	,
(	1331	)	,
(	1334	)	,
(	1337	)	,
(	1340	)	,
(	1343	)	,
(	1346	)	,
(	1349	)	,
(	1352	)	,
(	1355	)	,
(	1358	)	,
(	1361	)	,
(	1364	)	,
(	1367	)	,
(	1370	)	,
(	1373	)	,
(	1376	)	,
(	1379	)	,
(	1382	)	,
(	1385	)	,
(	1388	)	,
(	1391	)	,
(	1394	)	,
(	1398	)	,
(	1401	)	,
(	1404	)	,
(	1407	)	,
(	1410	)	,
(	1413	)	,
(	1416	)	,
(	1419	)	,
(	1422	)	,
(	1426	)	,
(	1429	)	,
(	1432	)	,
(	1435	)	,
(	1438	)	,
(	1441	)	,
(	1445	)	,
(	1448	)	,
(	1451	)	,
(	1454	)	,
(	1457	)	,
(	1461	)	,
(	1464	)	,
(	1467	)	,
(	1470	)	,
(	1473	)	,
(	1477	)	,
(	1480	)	,
(	1483	)	,
(	1487	)	,
(	1490	)	,
(	1493	)	,
(	1496	)	,
(	1500	)	,
(	1503	)	,
(	1506	)	,
(	1510	)	,
(	1513	)	,
(	1516	)	,
(	1520	)	,
(	1523	)	,
(	1526	)	,
(	1530	)	,
(	1533	)	,
(	1537	)	,
(	1540	)	,
(	1543	)	,
(	1547	)	,
(	1550	)	,
(	1554	)	,
(	1557	)	,
(	1560	)	,
(	1564	)	,
(	1567	)	,
(	1571	)	,
(	1574	)	,
(	1578	)	,
(	1581	)	,
(	1585	)	,
(	1588	)	,
(	1592	)	,
(	1595	)	,
(	1599	)	,
(	1602	)	,
(	1606	)	,
(	1609	)	,
(	1613	)	,
(	1616	)	,
(	1620	)	,
(	1624	)	,
(	1627	)	,
(	1631	)	,
(	1634	)	,
(	1638	)	,
(	1642	)	,
(	1645	)	,
(	1649	)	,
(	1652	)	,
(	1656	)	,
(	1660	)	,
(	1663	)	,
(	1667	)	,
(	1671	)	,
(	1674	)	,
(	1678	)	,
(	1682	)	,
(	1685	)	,
(	1689	)	,
(	1693	)	,
(	1697	)	,
(	1700	)	,
(	1704	)	,
(	1708	)	,
(	1712	)	,
(	1715	)	,
(	1719	)	,
(	1723	)	,
(	1727	)	,
(	1730	)	,
(	1734	)	,
(	1738	)	,
(	1742	)	,
(	1746	)	,
(	1750	)	,
(	1753	)	,
(	1757	)	,
(	1761	)	,
(	1765	)	,
(	1769	)	,
(	1773	)	,
(	1777	)	,
(	1781	)	,
(	1784	)	,
(	1788	)	,
(	1792	)	,
(	1796	)	,
(	1800	)	,
(	1804	)	,
(	1808	)	,
(	1812	)	,
(	1816	)	,
(	1820	)	,
(	1824	)	,
(	1828	)	,
(	1832	)	,
(	1836	)	,
(	1840	)	,
(	1844	)	,
(	1848	)	,
(	1852	)	,
(	1856	)	,
(	1860	)	,
(	1864	)	,
(	1868	)	,
(	1872	)	,
(	1877	)	,
(	1881	)	,
(	1885	)	,
(	1889	)	,
(	1893	)	,
(	1897	)	,
(	1901	)	,
(	1905	)	,
(	1910	)	,
(	1914	)	,
(	1918	)	,
(	1922	)	,
(	1926	)	,
(	1931	)	,
(	1935	)	,
(	1939	)	,
(	1943	)	,
(	1947	)	,
(	1952	)	,
(	1956	)	,
(	1960	)	,
(	1965	)	,
(	1969	)	,
(	1973	)	,
(	1977	)	,
(	1982	)	,
(	1986	)	,
(	1990	)	,
(	1995	)	,
(	1999	)	,
(	2003	)	,
(	2008	)	,
(	2012	)	,
(	2016	)	,
(	2021	)	,
(	2025	)	,
(	2030	)	,
(	2034	)	,
(	2038	)	,
(	2043	)	,
(	2047	)	,
(	2052	)	,
(	2056	)	,
(	2061	)	,
(	2065	)	,
(	2070	)	,
(	2074	)	,
(	2079	)	,
(	2083	)	,
(	2088	)	,
(	2092	)	,
(	2097	)	,
(	2101	)	,
(	2106	)	,
(	2110	)	,
(	2115	)	,
(	2120	)	,
(	2124	)	,
(	2129	)	,
(	2133	)	,
(	2138	)	,
(	2143	)	,
(	2147	)	,
(	2152	)	,
(	2156	)	,
(	2161	)	,
(	2166	)	,
(	2170	)	,
(	2175	)	,
(	2180	)	,
(	2185	)	,
(	2189	)	,
(	2194	)	,
(	2199	)	,
(	2203	)	,
(	2208	)	,
(	2213	)	,
(	2218	)	,
(	2222	)	,
(	2227	)	,
(	2232	)	,
(	2237	)	,
(	2242	)	,
(	2246	)	,
(	2251	)	,
(	2256	)	,
(	2261	)	,
(	2266	)	,
(	2271	)	,
(	2276	)	,
(	2280	)	,
(	2285	)	,
(	2290	)	,
(	2295	)	,
(	2300	)	,
(	2305	)	,
(	2310	)	,
(	2315	)	,
(	2320	)	,
(	2325	)	,
(	2330	)	,
(	2335	)	,
(	2340	)	,
(	2345	)	,
(	2350	)	,
(	2355	)	,
(	2360	)	,
(	2365	)	,
(	2370	)	,
(	2375	)	,
(	2380	)	,
(	2385	)	,
(	2390	)	,
(	2395	)	,
(	2401	)	,
(	2406	)	,
(	2411	)	,
(	2416	)	,
(	2421	)	,
(	2426	)	,
(	2431	)	,
(	2437	)	,
(	2442	)	,
(	2447	)	,
(	2452	)	,
(	2457	)	,
(	2463	)	,
(	2468	)	,
(	2473	)	,
(	2478	)	,
(	2484	)	,
(	2489	)	,
(	2494	)	,
(	2499	)	,
(	2505	)	,
(	2510	)	,
(	2515	)	,
(	2521	)	,
(	2526	)	,
(	2531	)	,
(	2537	)	,
(	2542	)	,
(	2548	)	,
(	2553	)	,
(	2558	)	,
(	2564	)	,
(	2569	)	,
(	2575	)	,
(	2580	)	,
(	2585	)	,
(	2591	)	,
(	2596	)	,
(	2602	)	,
(	2607	)	,
(	2613	)	,
(	2618	)	,
(	2624	)	,
(	2629	)	,
(	2635	)	,
(	2641	)	,
(	2646	)	,
(	2652	)	,
(	2657	)	,
(	2663	)	,
(	2668	)	,
(	2674	)	,
(	2680	)	,
(	2685	)	,
(	2691	)	,
(	2697	)	,
(	2702	)	,
(	2708	)	,
(	2714	)	,
(	2719	)	,
(	2725	)	,
(	2731	)	,
(	2736	)	,
(	2742	)	,
(	2748	)	,
(	2754	)	,
(	2759	)	,
(	2765	)	,
(	2771	)	,
(	2777	)	,
(	2783	)	,
(	2788	)	,
(	2794	)	,
(	2800	)	,
(	2806	)	,
(	2812	)	,
(	2818	)	,
(	2824	)	,
(	2829	)	,
(	2835	)	,
(	2841	)	,
(	2847	)	,
(	2853	)	,
(	2859	)	,
(	2865	)	,
(	2871	)	,
(	2877	)	,
(	2883	)	,
(	2889	)	,
(	2895	)	,
(	2901	)	,
(	2907	)	,
(	2913	)	,
(	2919	)	,
(	2925	)	,
(	2931	)	,
(	2937	)	,
(	2943	)	,
(	2949	)	,
(	2955	)	,
(	2962	)	,
(	2968	)	,
(	2974	)	,
(	2980	)	,
(	2986	)	,
(	2992	)	,
(	2999	)	,
(	3005	)	,
(	3011	)	,
(	3017	)	,
(	3023	)	,
(	3030	)	,
(	3036	)	,
(	3042	)	,
(	3048	)	,
(	3055	)	,
(	3061	)	,
(	3067	)	,
(	3074	)	,
(	3080	)	,
(	3086	)	,
(	3093	)	,
(	3099	)	,
(	3105	)	,
(	3112	)	,
(	3118	)	,
(	3125	)	,
(	3131	)	,
(	3137	)	,
(	3144	)	,
(	3150	)	,
(	3157	)	,
(	3163	)	,
(	3170	)	,
(	3176	)	,
(	3183	)	,
(	3189	)	,
(	3196	)	,
(	3202	)	,
(	3209	)	,
(	3215	)	,
(	3222	)	,
(	3228	)	,
(	3235	)	,
(	3242	)	,
(	3248	)	,
(	3255	)	,
(	3262	)	,
(	3268	)	,
(	3275	)	,
(	3281	)	,
(	3288	)	,
(	3295	)	,
(	3302	)	,
(	3308	)	,
(	3315	)	,
(	3322	)	,
(	3328	)	,
(	3335	)	,
(	3342	)	,
(	3349	)	,
(	3356	)	,
(	3362	)	,
(	3369	)	,
(	3376	)	,
(	3383	)	,
(	3390	)	,
(	3397	)	,
(	3403	)	,
(	3410	)	,
(	3417	)	,
(	3424	)	,
(	3431	)	,
(	3438	)	,
(	3445	)	,
(	3452	)	,
(	3459	)	,
(	3466	)	,
(	3473	)	,
(	3480	)	,
(	3487	)	,
(	3494	)	,
(	3501	)	,
(	3508	)	,
(	3515	)	,
(	3522	)	,
(	3529	)	,
(	3536	)	,
(	3543	)	,
(	3551	)	,
(	3558	)	,
(	3565	)	,
(	3572	)	,
(	3579	)	,
(	3586	)	,
(	3593	)	,
(	3601	)	,
(	3608	)	,
(	3615	)	,
(	3622	)	,
(	3630	)	,
(	3637	)	,
(	3644	)	,
(	3651	)	,
(	3659	)	,
(	3666	)	,
(	3673	)	,
(	3681	)	,
(	3688	)	,
(	3695	)	,
(	3703	)	,
(	3710	)	,
(	3718	)	,
(	3725	)	,
(	3732	)	,
(	3740	)	,
(	3747	)	,
(	3755	)	,
(	3762	)	,
(	3770	)	,
(	3777	)	,
(	3785	)	,
(	3792	)	,
(	3800	)	,
(	3807	)	,
(	3815	)	,
(	3822	)	,
(	3830	)	,
(	3837	)	,
(	3845	)	,
(	3853	)	,
(	3860	)	,
(	3868	)	,
(	3876	)	,
(	3883	)	,
(	3891	)	,
(	3899	)	,
(	3906	)	,
(	3914	)	,
(	3922	)	,
(	3930	)	,
(	3937	)	,
(	3945	)	,
(	3953	)	,
(	3961	)	,
(	3968	)	,
(	3976	)	,
(	3984	)	,
(	3992	)	,
(	4000	)	,
(	4008	)	,
(	4015	)	,
(	4023	)	,
(	4031	)	,
(	4039	)	,
(	4047	)	,
(	4055	)	,
(	4063	)	,
(	4071	)	,
(	4079	)	,
(	4087	)	,
(	4095	)	,
(	4103	)	,
(	4111	)	,
(	4119	)	,
(	4127	)	,
(	4135	)	,
(	4143	)	,
(	4151	)	,
(	4159	)	,
(	4167	)	,
(	4176	)	,
(	4184	)	,
(	4192	)	,
(	4200	)	,
(	4208	)	,
(	4216	)	,
(	4225	)	,
(	4233	)	,
(	4241	)	,
(	4249	)	,
(	4258	)	,
(	4266	)	,
(	4274	)	,
(	4282	)	,
(	4291	)	,
(	4299	)	,
(	4307	)	,
(	4316	)	,
(	4324	)	,
(	4332	)	,
(	4341	)	,
(	4349	)	,
(	4358	)	,
(	4366	)	,
(	4374	)	,
(	4383	)	,
(	4391	)	,
(	4400	)	,
(	4408	)	,
(	4417	)	,
(	4425	)	,
(	4434	)	,
(	4442	)	,
(	4451	)	,
(	4460	)	,
(	4468	)	,
(	4477	)	,
(	4485	)	,
(	4494	)	,
(	4503	)	,
(	4511	)	,
(	4520	)	,
(	4529	)	,
(	4537	)	,
(	4546	)	,
(	4555	)	,
(	4563	)	,
(	4572	)	,
(	4581	)	,
(	4590	)	,
(	4598	)	,
(	4607	)	,
(	4616	)	,
(	4625	)	,
(	4634	)	,
(	4643	)	,
(	4651	)	,
(	4660	)	,
(	4669	)	,
(	4678	)	,
(	4687	)	,
(	4696	)	,
(	4705	)	,
(	4714	)	,
(	4723	)	,
(	4732	)	,
(	4741	)	,
(	4750	)	,
(	4759	)	,
(	4768	)	,
(	4777	)	,
(	4786	)	,
(	4795	)	,
(	4804	)	,
(	4813	)	,
(	4823	)	,
(	4832	)	,
(	4841	)	,
(	4850	)	,
(	4859	)	,
(	4868	)	,
(	4878	)	,
(	4887	)	,
(	4896	)	,
(	4905	)	,
(	4915	)	,
(	4924	)	,
(	4933	)	,
(	4942	)	,
(	4952	)	,
(	4961	)	,
(	4970	)	,
(	4980	)	,
(	4989	)	,
(	4999	)	,
(	5008	)	,
(	5017	)	,
(	5027	)	,
(	5036	)	,
(	5046	)	,
(	5055	)	,
(	5065	)	,
(	5074	)	,
(	5084	)	,
(	5093	)	,
(	5103	)	,
(	5112	)	,
(	5122	)	,
(	5131	)	,
(	5141	)	,
(	5151	)	,
(	5160	)	,
(	5170	)	,
(	5180	)	,
(	5189	)	,
(	5199	)	,
(	5209	)	,
(	5218	)	,
(	5228	)	,
(	5238	)	,
(	5248	)	,
(	5257	)	,
(	5267	)	,
(	5277	)	,
(	5287	)	,
(	5297	)	,
(	5307	)	,
(	5316	)	,
(	5326	)	,
(	5336	)	,
(	5346	)	,
(	5356	)	,
(	5366	)	,
(	5376	)	,
(	5386	)	,
(	5396	)	,
(	5406	)	,
(	5416	)	,
(	5426	)	,
(	5436	)	,
(	5446	)	,
(	5456	)	,
(	5466	)	,
(	5476	)	,
(	5486	)	,
(	5496	)	,
(	5507	)	,
(	5517	)	,
(	5527	)	,
(	5537	)	,
(	5547	)	,
(	5557	)	,
(	5568	)	,
(	5578	)	,
(	5588	)	,
(	5598	)	,
(	5609	)	,
(	5619	)	,
(	5629	)	,
(	5640	)	,
(	5650	)	,
(	5660	)	,
(	5671	)	,
(	5681	)	,
(	5692	)	,
(	5702	)	,
(	5712	)	,
(	5723	)	,
(	5733	)	,
(	5744	)	,
(	5754	)	,
(	5765	)	,
(	5775	)	,
(	5786	)	,
(	5797	)	,
(	5807	)	,
(	5818	)	,
(	5828	)	,
(	5839	)	,
(	5850	)	,
(	5860	)	,
(	5871	)	,
(	5882	)	,
(	5892	)	,
(	5903	)	,
(	5914	)	,
(	5924	)	,
(	5935	)	,
(	5946	)	,
(	5957	)	,
(	5968	)	,
(	5978	)	,
(	5989	)	,
(	6000	)	,
(	6011	)	,
(	6022	)	,
(	6033	)	,
(	6044	)	,
(	6055	)	,
(	6066	)	,
(	6076	)	,
(	6087	)	,
(	6098	)	,
(	6109	)	,
(	6120	)	,
(	6132	)	,
(	6143	)	,
(	6154	)		-- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 6154 (61.54 cm)

);


end package LUT_pkg;
