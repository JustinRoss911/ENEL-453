library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_flashing_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant d2freq_LUT : array_1d := (

(	65152	)	,
(	65138	)	,
(	65124	)	,
(	65111	)	,
(	65097	)	,
(	65083	)	,
(	65069	)	,
(	65055	)	,
(	65042	)	,
(	65028	)	,
(	65014	)	,
(	65000	)	,
(	64987	)	,
(	64973	)	,
(	64959	)	,
(	64945	)	,
(	64931	)	,
(	64918	)	,
(	64904	)	,
(	64890	)	,
(	64876	)	,
(	64862	)	,
(	64849	)	,
(	64835	)	,
(	64821	)	,
(	64807	)	,
(	64793	)	,
(	64780	)	,
(	64766	)	,
(	64752	)	,
(	64738	)	,
(	64725	)	,
(	64711	)	,
(	64697	)	,
(	64683	)	,
(	64669	)	,
(	64656	)	,
(	64642	)	,
(	64628	)	,
(	64614	)	,
(	64600	)	,
(	64587	)	,
(	64573	)	,
(	64559	)	,
(	64545	)	,
(	64531	)	,
(	64518	)	,
(	64504	)	,
(	64490	)	,
(	64476	)	,
(	64463	)	,
(	64449	)	,
(	64435	)	,
(	64421	)	,
(	64407	)	,
(	64394	)	,
(	64380	)	,
(	64366	)	,
(	64352	)	,
(	64338	)	,
(	64325	)	,
(	64311	)	,
(	64297	)	,
(	64283	)	,
(	64270	)	,
(	64256	)	,
(	64242	)	,
(	64228	)	,
(	64214	)	,
(	64201	)	,
(	64187	)	,
(	64173	)	,
(	64159	)	,
(	64145	)	,
(	64132	)	,
(	64118	)	,
(	64104	)	,
(	64090	)	,
(	64076	)	,
(	64063	)	,
(	64049	)	,
(	64035	)	,
(	64021	)	,
(	64008	)	,
(	63994	)	,
(	63980	)	,
(	63966	)	,
(	63952	)	,
(	63939	)	,
(	63925	)	,
(	63911	)	,
(	63897	)	,
(	63883	)	,
(	63870	)	,
(	63856	)	,
(	63842	)	,
(	63828	)	,
(	63814	)	,
(	63801	)	,
(	63787	)	,
(	63773	)	,
(	63759	)	,
(	63746	)	,
(	63732	)	,
(	63718	)	,
(	63704	)	,
(	63690	)	,
(	63677	)	,
(	63663	)	,
(	63649	)	,
(	63635	)	,
(	63621	)	,
(	63608	)	,
(	63594	)	,
(	63580	)	,
(	63566	)	,
(	63552	)	,
(	63539	)	,
(	63525	)	,
(	63511	)	,
(	63497	)	,
(	63484	)	,
(	63470	)	,
(	63456	)	,
(	63442	)	,
(	63428	)	,
(	63415	)	,
(	63401	)	,
(	63387	)	,
(	63373	)	,
(	63359	)	,
(	63346	)	,
(	63332	)	,
(	63318	)	,
(	63304	)	,
(	63290	)	,
(	63277	)	,
(	63263	)	,
(	63249	)	,
(	63235	)	,
(	63222	)	,
(	63208	)	,
(	63194	)	,
(	63180	)	,
(	63166	)	,
(	63153	)	,
(	63139	)	,
(	63125	)	,
(	63111	)	,
(	63097	)	,
(	63084	)	,
(	63070	)	,
(	63056	)	,
(	63042	)	,
(	63028	)	,
(	63015	)	,
(	63001	)	,
(	62987	)	,
(	62973	)	,
(	62960	)	,
(	62946	)	,
(	62932	)	,
(	62918	)	,
(	62904	)	,
(	62891	)	,
(	62877	)	,
(	62863	)	,
(	62849	)	,
(	62835	)	,
(	62822	)	,
(	62808	)	,
(	62794	)	,
(	62780	)	,
(	62767	)	,
(	62753	)	,
(	62739	)	,
(	62725	)	,
(	62711	)	,
(	62698	)	,
(	62684	)	,
(	62670	)	,
(	62656	)	,
(	62642	)	,
(	62629	)	,
(	62615	)	,
(	62601	)	,
(	62587	)	,
(	62573	)	,
(	62560	)	,
(	62546	)	,
(	62532	)	,
(	62518	)	,
(	62505	)	,
(	62491	)	,
(	62477	)	,
(	62463	)	,
(	62449	)	,
(	62436	)	,
(	62422	)	,
(	62408	)	,
(	62394	)	,
(	62380	)	,
(	62367	)	,
(	62353	)	,
(	62339	)	,
(	62325	)	,
(	62311	)	,
(	62298	)	,
(	62284	)	,
(	62270	)	,
(	62256	)	,
(	62243	)	,
(	62229	)	,
(	62215	)	,
(	62201	)	,
(	62187	)	,
(	62174	)	,
(	62160	)	,
(	62146	)	,
(	62132	)	,
(	62118	)	,
(	62105	)	,
(	62091	)	,
(	62077	)	,
(	62063	)	,
(	62049	)	,
(	62036	)	,
(	62022	)	,
(	62008	)	,
(	61994	)	,
(	61981	)	,
(	61967	)	,
(	61953	)	,
(	61939	)	,
(	61925	)	,
(	61912	)	,
(	61898	)	,
(	61884	)	,
(	61870	)	,
(	61856	)	,
(	61843	)	,
(	61829	)	,
(	61815	)	,
(	61801	)	,
(	61787	)	,
(	61774	)	,
(	61760	)	,
(	61746	)	,
(	61732	)	,
(	61719	)	,
(	61705	)	,
(	61691	)	,
(	61677	)	,
(	61663	)	,
(	61650	)	,
(	61636	)	,
(	61622	)	,
(	61608	)	,
(	61594	)	,
(	61581	)	,
(	61567	)	,
(	61553	)	,
(	61539	)	,
(	61525	)	,
(	61512	)	,
(	61498	)	,
(	61484	)	,
(	61470	)	,
(	61457	)	,
(	61443	)	,
(	61429	)	,
(	61415	)	,
(	61401	)	,
(	61388	)	,
(	61374	)	,
(	61360	)	,
(	61346	)	,
(	61332	)	,
(	61319	)	,
(	61305	)	,
(	61291	)	,
(	61277	)	,
(	61264	)	,
(	61250	)	,
(	61236	)	,
(	61222	)	,
(	61208	)	,
(	61195	)	,
(	61181	)	,
(	61167	)	,
(	61153	)	,
(	61139	)	,
(	61126	)	,
(	61112	)	,
(	61098	)	,
(	61084	)	,
(	61070	)	,
(	61057	)	,
(	61043	)	,
(	61029	)	,
(	61015	)	,
(	61002	)	,
(	60988	)	,
(	60974	)	,
(	60960	)	,
(	60946	)	,
(	60933	)	,
(	60919	)	,
(	60905	)	,
(	60891	)	,
(	60877	)	,
(	60864	)	,
(	60850	)	,
(	60836	)	,
(	60822	)	,
(	60808	)	,
(	60795	)	,
(	60781	)	,
(	60767	)	,
(	60753	)	,
(	60740	)	,
(	60726	)	,
(	60712	)	,
(	60698	)	,
(	60684	)	,
(	60671	)	,
(	60657	)	,
(	60643	)	,
(	60629	)	,
(	60615	)	,
(	60602	)	,
(	60588	)	,
(	60574	)	,
(	60560	)	,
(	60546	)	,
(	60533	)	,
(	60519	)	,
(	60505	)	,
(	60491	)	,
(	60478	)	,
(	60464	)	,
(	60450	)	,
(	60436	)	,
(	60422	)	,
(	60409	)	,
(	60395	)	,
(	60381	)	,
(	60367	)	,
(	60353	)	,
(	60340	)	,
(	60326	)	,
(	60312	)	,
(	60298	)	,
(	60284	)	,
(	60271	)	,
(	60257	)	,
(	60243	)	,
(	60229	)	,
(	60216	)	,
(	60202	)	,
(	60188	)	,
(	60174	)	,
(	60160	)	,
(	60147	)	,
(	60133	)	,
(	60119	)	,
(	60105	)	,
(	60091	)	,
(	60078	)	,
(	60064	)	,
(	60050	)	,
(	60036	)	,
(	60022	)	,
(	60009	)	,
(	59995	)	,
(	59981	)	,
(	59967	)	,
(	59954	)	,
(	59940	)	,
(	59926	)	,
(	59912	)	,
(	59898	)	,
(	59885	)	,
(	59871	)	,
(	59857	)	,
(	59843	)	,
(	59829	)	,
(	59816	)	,
(	59802	)	,
(	59788	)	,
(	59774	)	,
(	59761	)	,
(	59747	)	,
(	59733	)	,
(	59719	)	,
(	59705	)	,
(	59692	)	,
(	59678	)	,
(	59664	)	,
(	59650	)	,
(	59636	)	,
(	59623	)	,
(	59609	)	,
(	59595	)	,
(	59581	)	,
(	59567	)	,
(	59554	)	,
(	59540	)	,
(	59526	)	,
(	59512	)	,
(	59499	)	,
(	59485	)	,
(	59471	)	,
(	59457	)	,
(	59443	)	,
(	59430	)	,
(	59416	)	,
(	59402	)	,
(	59388	)	,
(	59374	)	,
(	59361	)	,
(	59347	)	,
(	59333	)	,
(	59319	)	,
(	59305	)	,
(	59292	)	,
(	59278	)	,
(	59264	)	,
(	59250	)	,
(	59237	)	,
(	59223	)	,
(	59209	)	,
(	59195	)	,
(	59181	)	,
(	59168	)	,
(	59154	)	,
(	59140	)	,
(	59126	)	,
(	59112	)	,
(	59099	)	,
(	59085	)	,
(	59071	)	,
(	59057	)	,
(	59043	)	,
(	59030	)	,
(	59016	)	,
(	59002	)	,
(	58988	)	,
(	58975	)	,
(	58961	)	,
(	58947	)	,
(	58933	)	,
(	58919	)	,
(	58906	)	,
(	58892	)	,
(	58878	)	,
(	58864	)	,
(	58850	)	,
(	58837	)	,
(	58823	)	,
(	58809	)	,
(	58795	)	,
(	58781	)	,
(	58768	)	,
(	58754	)	,
(	58740	)	,
(	58726	)	,
(	58713	)	,
(	58699	)	,
(	58685	)	,
(	58671	)	,
(	58657	)	,
(	58644	)	,
(	58630	)	,
(	58616	)	,
(	58602	)	,
(	58588	)	,
(	58575	)	,
(	58561	)	,
(	58547	)	,
(	58533	)	,
(	58519	)	,
(	58506	)	,
(	58492	)	,
(	58478	)	,
(	58464	)	,
(	58451	)	,
(	58437	)	,
(	58423	)	,
(	58409	)	,
(	58395	)	,
(	58382	)	,
(	58368	)	,
(	58354	)	,
(	58340	)	,
(	58326	)	,
(	58313	)	,
(	58299	)	,
(	58285	)	,
(	58271	)	,
(	58258	)	,
(	58244	)	,
(	58230	)	,
(	58216	)	,
(	58202	)	,
(	58189	)	,
(	58175	)	,
(	58161	)	,
(	58147	)	,
(	58133	)	,
(	58120	)	,
(	58106	)	,
(	58092	)	,
(	58078	)	,
(	58064	)	,
(	58051	)	,
(	58037	)	,
(	58023	)	,
(	58009	)	,
(	57996	)	,
(	57982	)	,
(	57968	)	,
(	57954	)	,
(	57940	)	,
(	57927	)	,
(	57913	)	,
(	57899	)	,
(	57885	)	,
(	57871	)	,
(	57858	)	,
(	57844	)	,
(	57830	)	,
(	57816	)	,
(	57802	)	,
(	57789	)	,
(	57775	)	,
(	57761	)	,
(	57747	)	,
(	57734	)	,
(	57720	)	,
(	57706	)	,
(	57692	)	,
(	57678	)	,
(	57665	)	,
(	57651	)	,
(	57637	)	,
(	57623	)	,
(	57609	)	,
(	57596	)	,
(	57582	)	,
(	57568	)	,
(	57554	)	,
(	57540	)	,
(	57527	)	,
(	57513	)	,
(	57499	)	,
(	57485	)	,
(	57472	)	,
(	57458	)	,
(	57444	)	,
(	57430	)	,
(	57416	)	,
(	57403	)	,
(	57389	)	,
(	57375	)	,
(	57361	)	,
(	57347	)	,
(	57334	)	,
(	57320	)	,
(	57306	)	,
(	57292	)	,
(	57278	)	,
(	57265	)	,
(	57251	)	,
(	57237	)	,
(	57223	)	,
(	57210	)	,
(	57196	)	,
(	57182	)	,
(	57168	)	,
(	57154	)	,
(	57141	)	,
(	57127	)	,
(	57113	)	,
(	57099	)	,
(	57085	)	,
(	57072	)	,
(	57058	)	,
(	57044	)	,
(	57030	)	,
(	57016	)	,
(	57003	)	,
(	56989	)	,
(	56975	)	,
(	56961	)	,
(	56948	)	,
(	56934	)	,
(	56920	)	,
(	56906	)	,
(	56892	)	,
(	56879	)	,
(	56865	)	,
(	56851	)	,
(	56837	)	,
(	56823	)	,
(	56810	)	,
(	56796	)	,
(	56782	)	,
(	56768	)	,
(	56754	)	,
(	56741	)	,
(	56727	)	,
(	56713	)	,
(	56699	)	,
(	56686	)	,
(	56672	)	,
(	56658	)	,
(	56644	)	,
(	56630	)	,
(	56617	)	,
(	56603	)	,
(	56589	)	,
(	56575	)	,
(	56561	)	,
(	56548	)	,
(	56534	)	,
(	56520	)	,
(	56506	)	,
(	56493	)	,
(	56479	)	,
(	56465	)	,
(	56451	)	,
(	56437	)	,
(	56424	)	,
(	56410	)	,
(	56396	)	,
(	56382	)	,
(	56368	)	,
(	56355	)	,
(	56341	)	,
(	56327	)	,
(	56313	)	,
(	56299	)	,
(	56286	)	,
(	56272	)	,
(	56258	)	,
(	56244	)	,
(	56231	)	,
(	56217	)	,
(	56203	)	,
(	56189	)	,
(	56175	)	,
(	56162	)	,
(	56148	)	,
(	56134	)	,
(	56120	)	,
(	56106	)	,
(	56093	)	,
(	56079	)	,
(	56065	)	,
(	56051	)	,
(	56037	)	,
(	56024	)	,
(	56010	)	,
(	55996	)	,
(	55982	)	,
(	55969	)	,
(	55955	)	,
(	55941	)	,
(	55927	)	,
(	55913	)	,
(	55900	)	,
(	55886	)	,
(	55872	)	,
(	55858	)	,
(	55844	)	,
(	55831	)	,
(	55817	)	,
(	55803	)	,
(	55789	)	,
(	55775	)	,
(	55762	)	,
(	55748	)	,
(	55734	)	,
(	55720	)	,
(	55707	)	,
(	55693	)	,
(	55679	)	,
(	55665	)	,
(	55651	)	,
(	55638	)	,
(	55624	)	,
(	55610	)	,
(	55596	)	,
(	55582	)	,
(	55569	)	,
(	55555	)	,
(	55541	)	,
(	55527	)	,
(	55513	)	,
(	55500	)	,
(	55486	)	,
(	55472	)	,
(	55458	)	,
(	55445	)	,
(	55431	)	,
(	55417	)	,
(	55403	)	,
(	55389	)	,
(	55376	)	,
(	55362	)	,
(	55348	)	,
(	55334	)	,
(	55320	)	,
(	55307	)	,
(	55293	)	,
(	55279	)	,
(	55265	)	,
(	55251	)	,
(	55238	)	,
(	55224	)	,
(	55210	)	,
(	55196	)	,
(	55183	)	,
(	55169	)	,
(	55155	)	,
(	55141	)	,
(	55127	)	,
(	55114	)	,
(	55100	)	,
(	55086	)	,
(	55072	)	,
(	55058	)	,
(	55045	)	,
(	55031	)	,
(	55017	)	,
(	55003	)	,
(	54990	)	,
(	54976	)	,
(	54962	)	,
(	54948	)	,
(	54934	)	,
(	54921	)	,
(	54907	)	,
(	54893	)	,
(	54879	)	,
(	54865	)	,
(	54852	)	,
(	54838	)	,
(	54824	)	,
(	54810	)	,
(	54796	)	,
(	54783	)	,
(	54769	)	,
(	54755	)	,
(	54741	)	,
(	54728	)	,
(	54714	)	,
(	54700	)	,
(	54686	)	,
(	54672	)	,
(	54659	)	,
(	54645	)	,
(	54631	)	,
(	54617	)	,
(	54603	)	,
(	54590	)	,
(	54576	)	,
(	54562	)	,
(	54548	)	,
(	54534	)	,
(	54521	)	,
(	54507	)	,
(	54493	)	,
(	54479	)	,
(	54466	)	,
(	54452	)	,
(	54438	)	,
(	54424	)	,
(	54410	)	,
(	54397	)	,
(	54383	)	,
(	54369	)	,
(	54355	)	,
(	54341	)	,
(	54328	)	,
(	54314	)	,
(	54300	)	,
(	54286	)	,
(	54272	)	,
(	54259	)	,
(	54245	)	,
(	54231	)	,
(	54217	)	,
(	54204	)	,
(	54190	)	,
(	54176	)	,
(	54162	)	,
(	54148	)	,
(	54135	)	,
(	54121	)	,
(	54107	)	,
(	54093	)	,
(	54079	)	,
(	54066	)	,
(	54052	)	,
(	54038	)	,
(	54024	)	,
(	54010	)	,
(	53997	)	,
(	53983	)	,
(	53969	)	,
(	53955	)	,
(	53942	)	,
(	53928	)	,
(	53914	)	,
(	53900	)	,
(	53886	)	,
(	53873	)	,
(	53859	)	,
(	53845	)	,
(	53831	)	,
(	53817	)	,
(	53804	)	,
(	53790	)	,
(	53776	)	,
(	53762	)	,
(	53748	)	,
(	53735	)	,
(	53721	)	,
(	53707	)	,
(	53693	)	,
(	53680	)	,
(	53666	)	,
(	53652	)	,
(	53638	)	,
(	53624	)	,
(	53611	)	,
(	53597	)	,
(	53583	)	,
(	53569	)	,
(	53555	)	,
(	53542	)	,
(	53528	)	,
(	53514	)	,
(	53500	)	,
(	53487	)	,
(	53473	)	,
(	53459	)	,
(	53445	)	,
(	53431	)	,
(	53418	)	,
(	53404	)	,
(	53390	)	,
(	53376	)	,
(	53362	)	,
(	53349	)	,
(	53335	)	,
(	53321	)	,
(	53307	)	,
(	53293	)	,
(	53280	)	,
(	53266	)	,
(	53252	)	,
(	53238	)	,
(	53225	)	,
(	53211	)	,
(	53197	)	,
(	53183	)	,
(	53169	)	,
(	53156	)	,
(	53142	)	,
(	53128	)	,
(	53114	)	,
(	53100	)	,
(	53087	)	,
(	53073	)	,
(	53059	)	,
(	53045	)	,
(	53031	)	,
(	53018	)	,
(	53004	)	,
(	52990	)	,
(	52976	)	,
(	52963	)	,
(	52949	)	,
(	52935	)	,
(	52921	)	,
(	52907	)	,
(	52894	)	,
(	52880	)	,
(	52866	)	,
(	52852	)	,
(	52838	)	,
(	52825	)	,
(	52811	)	,
(	52797	)	,
(	52783	)	,
(	52769	)	,
(	52756	)	,
(	52742	)	,
(	52728	)	,
(	52714	)	,
(	52701	)	,
(	52687	)	,
(	52673	)	,
(	52659	)	,
(	52645	)	,
(	52632	)	,
(	52618	)	,
(	52604	)	,
(	52590	)	,
(	52576	)	,
(	52563	)	,
(	52549	)	,
(	52535	)	,
(	52521	)	,
(	52507	)	,
(	52494	)	,
(	52480	)	,
(	52466	)	,
(	52452	)	,
(	52439	)	,
(	52425	)	,
(	52411	)	,
(	52397	)	,
(	52383	)	,
(	52370	)	,
(	52356	)	,
(	52342	)	,
(	52328	)	,
(	52314	)	,
(	52301	)	,
(	52287	)	,
(	52273	)	,
(	52259	)	,
(	52245	)	,
(	52232	)	,
(	52218	)	,
(	52204	)	,
(	52190	)	,
(	52177	)	,
(	52163	)	,
(	52149	)	,
(	52135	)	,
(	52121	)	,
(	52108	)	,
(	52094	)	,
(	52080	)	,
(	52066	)	,
(	52052	)	,
(	52039	)	,
(	52025	)	,
(	52011	)	,
(	51997	)	,
(	51984	)	,
(	51970	)	,
(	51956	)	,
(	51942	)	,
(	51928	)	,
(	51915	)	,
(	51901	)	,
(	51887	)	,
(	51873	)	,
(	51859	)	,
(	51846	)	,
(	51832	)	,
(	51818	)	,
(	51804	)	,
(	51790	)	,
(	51777	)	,
(	51763	)	,
(	51749	)	,
(	51735	)	,
(	51722	)	,
(	51708	)	,
(	51694	)	,
(	51680	)	,
(	51666	)	,
(	51653	)	,
(	51639	)	,
(	51625	)	,
(	51611	)	,
(	51597	)	,
(	51584	)	,
(	51570	)	,
(	51556	)	,
(	51542	)	,
(	51528	)	,
(	51515	)	,
(	51501	)	,
(	51487	)	,
(	51473	)	,
(	51460	)	,
(	51446	)	,
(	51432	)	,
(	51418	)	,
(	51404	)	,
(	51391	)	,
(	51377	)	,
(	51363	)	,
(	51349	)	,
(	51335	)	,
(	51322	)	,
(	51308	)	,
(	51294	)	,
(	51280	)	,
(	51266	)	,
(	51253	)	,
(	51239	)	,
(	51225	)	,
(	51211	)	,
(	51198	)	,
(	51184	)	,
(	51170	)	,
(	51156	)	,
(	51142	)	,
(	51129	)	,
(	51115	)	,
(	51101	)	,
(	51087	)	,
(	51073	)	,
(	51060	)	,
(	51046	)	,
(	51032	)	,
(	51018	)	,
(	51004	)	,
(	50991	)	,
(	50977	)	,
(	50963	)	,
(	50949	)	,
(	50936	)	,
(	50922	)	,
(	50908	)	,
(	50894	)	,
(	50880	)	,
(	50867	)	,
(	50853	)	,
(	50839	)	,
(	50825	)	,
(	50811	)	,
(	50798	)	,
(	50784	)	,
(	50770	)	,
(	50756	)	,
(	50742	)	,
(	50729	)	,
(	50715	)	,
(	50701	)	,
(	50687	)	,
(	50674	)	,
(	50660	)	,
(	50646	)	,
(	50632	)	,
(	50618	)	,
(	50605	)	,
(	50591	)	,
(	50577	)	,
(	50563	)	,
(	50549	)	,
(	50536	)	,
(	50522	)	,
(	50508	)	,
(	50494	)	,
(	50481	)	,
(	50467	)	,
(	50453	)	,
(	50439	)	,
(	50425	)	,
(	50412	)	,
(	50398	)	,
(	50384	)	,
(	50370	)	,
(	50356	)	,
(	50343	)	,
(	50329	)	,
(	50315	)	,
(	50301	)	,
(	50287	)	,
(	50274	)	,
(	50260	)	,
(	50246	)	,
(	50232	)	,
(	50219	)	,
(	50205	)	,
(	50191	)	,
(	50177	)	,
(	50163	)	,
(	50150	)	,
(	50136	)	,
(	50122	)	,
(	50108	)	,
(	50094	)	,
(	50081	)	,
(	50067	)	,
(	50053	)	,
(	50039	)	,
(	50025	)	,
(	50012	)	,
(	49998	)	,
(	49984	)	,
(	49970	)	,
(	49957	)	,
(	49943	)	,
(	49929	)	,
(	49915	)	,
(	49901	)	,
(	49888	)	,
(	49874	)	,
(	49860	)	,
(	49846	)	,
(	49832	)	,
(	49819	)	,
(	49805	)	,
(	49791	)	,
(	49777	)	,
(	49763	)	,
(	49750	)	,
(	49736	)	,
(	49722	)	,
(	49708	)	,
(	49695	)	,
(	49681	)	,
(	49667	)	,
(	49653	)	,
(	49639	)	,
(	49626	)	,
(	49612	)	,
(	49598	)	,
(	49584	)	,
(	49570	)	,
(	49557	)	,
(	49543	)	,
(	49529	)	,
(	49515	)	,
(	49501	)	,
(	49488	)	,
(	49474	)	,
(	49460	)	,
(	49446	)	,
(	49433	)	,
(	49419	)	,
(	49405	)	,
(	49391	)	,
(	49377	)	,
(	49364	)	,
(	49350	)	,
(	49336	)	,
(	49322	)	,
(	49308	)	,
(	49295	)	,
(	49281	)	,
(	49267	)	,
(	49253	)	,
(	49239	)	,
(	49226	)	,
(	49212	)	,
(	49198	)	,
(	49184	)	,
(	49171	)	,
(	49157	)	,
(	49143	)	,
(	49129	)	,
(	49115	)	,
(	49102	)	,
(	49088	)	,
(	49074	)	,
(	49060	)	,
(	49046	)	,
(	49033	)	,
(	49019	)	,
(	49005	)	,
(	48991	)	,
(	48978	)	,
(	48964	)	,
(	48950	)	,
(	48936	)	,
(	48922	)	,
(	48909	)	,
(	48895	)	,
(	48881	)	,
(	48867	)	,
(	48853	)	,
(	48840	)	,
(	48826	)	,
(	48812	)	,
(	48798	)	,
(	48784	)	,
(	48771	)	,
(	48757	)	,
(	48743	)	,
(	48729	)	,
(	48716	)	,
(	48702	)	,
(	48688	)	,
(	48674	)	,
(	48660	)	,
(	48647	)	,
(	48633	)	,
(	48619	)	,
(	48605	)	,
(	48591	)	,
(	48578	)	,
(	48564	)	,
(	48550	)	,
(	48536	)	,
(	48522	)	,
(	48509	)	,
(	48495	)	,
(	48481	)	,
(	48467	)	,
(	48454	)	,
(	48440	)	,
(	48426	)	,
(	48412	)	,
(	48398	)	,
(	48385	)	,
(	48371	)	,
(	48357	)	,
(	48343	)	,
(	48329	)	,
(	48316	)	,
(	48302	)	,
(	48288	)	,
(	48274	)	,
(	48260	)	,
(	48247	)	,
(	48233	)	,
(	48219	)	,
(	48205	)	,
(	48192	)	,
(	48178	)	,
(	48164	)	,
(	48150	)	,
(	48136	)	,
(	48123	)	,
(	48109	)	,
(	48095	)	,
(	48081	)	,
(	48067	)	,
(	48054	)	,
(	48040	)	,
(	48026	)	,
(	48012	)	,
(	47998	)	,
(	47985	)	,
(	47971	)	,
(	47957	)	,
(	47943	)	,
(	47930	)	,
(	47916	)	,
(	47902	)	,
(	47888	)	,
(	47874	)	,
(	47861	)	,
(	47847	)	,
(	47833	)	,
(	47819	)	,
(	47805	)	,
(	47792	)	,
(	47778	)	,
(	47764	)	,
(	47750	)	,
(	47736	)	,
(	47723	)	,
(	47709	)	,
(	47695	)	,
(	47681	)	,
(	47668	)	,
(	47654	)	,
(	47640	)	,
(	47626	)	,
(	47612	)	,
(	47599	)	,
(	47585	)	,
(	47571	)	,
(	47557	)	,
(	47543	)	,
(	47530	)	,
(	47516	)	,
(	47502	)	,
(	47488	)	,
(	47475	)	,
(	47461	)	,
(	47447	)	,
(	47433	)	,
(	47419	)	,
(	47406	)	,
(	47392	)	,
(	47378	)	,
(	47364	)	,
(	47350	)	,
(	47337	)	,
(	47323	)	,
(	47309	)	,
(	47295	)	,
(	47281	)	,
(	47268	)	,
(	47254	)	,
(	47240	)	,
(	47226	)	,
(	47213	)	,
(	47199	)	,
(	47185	)	,
(	47171	)	,
(	47157	)	,
(	47144	)	,
(	47130	)	,
(	47116	)	,
(	47102	)	,
(	47088	)	,
(	47075	)	,
(	47061	)	,
(	47047	)	,
(	47033	)	,
(	47019	)	,
(	47006	)	,
(	46992	)	,
(	46978	)	,
(	46964	)	,
(	46951	)	,
(	46937	)	,
(	46923	)	,
(	46909	)	,
(	46895	)	,
(	46882	)	,
(	46868	)	,
(	46854	)	,
(	46840	)	,
(	46826	)	,
(	46813	)	,
(	46799	)	,
(	46785	)	,
(	46771	)	,
(	46757	)	,
(	46744	)	,
(	46730	)	,
(	46716	)	,
(	46702	)	,
(	46689	)	,
(	46675	)	,
(	46661	)	,
(	46647	)	,
(	46633	)	,
(	46620	)	,
(	46606	)	,
(	46592	)	,
(	46578	)	,
(	46564	)	,
(	46551	)	,
(	46537	)	,
(	46523	)	,
(	46509	)	,
(	46495	)	,
(	46482	)	,
(	46468	)	,
(	46454	)	,
(	46440	)	,
(	46427	)	,
(	46413	)	,
(	46399	)	,
(	46385	)	,
(	46371	)	,
(	46358	)	,
(	46344	)	,
(	46330	)	,
(	46316	)	,
(	46302	)	,
(	46289	)	,
(	46275	)	,
(	46261	)	,
(	46247	)	,
(	46233	)	,
(	46220	)	,
(	46206	)	,
(	46192	)	,
(	46178	)	,
(	46165	)	,
(	46151	)	,
(	46137	)	,
(	46123	)	,
(	46109	)	,
(	46096	)	,
(	46082	)	,
(	46068	)	,
(	46054	)	,
(	46040	)	,
(	46027	)	,
(	46013	)	,
(	45999	)	,
(	45985	)	,
(	45972	)	,
(	45958	)	,
(	45944	)	,
(	45930	)	,
(	45916	)	,
(	45903	)	,
(	45889	)	,
(	45875	)	,
(	45861	)	,
(	45847	)	,
(	45834	)	,
(	45820	)	,
(	45806	)	,
(	45792	)	,
(	45778	)	,
(	45765	)	,
(	45751	)	,
(	45737	)	,
(	45723	)	,
(	45710	)	,
(	45696	)	,
(	45682	)	,
(	45668	)	,
(	45654	)	,
(	45641	)	,
(	45627	)	,
(	45613	)	,
(	45599	)	,
(	45585	)	,
(	45572	)	,
(	45558	)	,
(	45544	)	,
(	45530	)	,
(	45516	)	,
(	45503	)	,
(	45489	)	,
(	45475	)	,
(	45461	)	,
(	45448	)	,
(	45434	)	,
(	45420	)	,
(	45406	)	,
(	45392	)	,
(	45379	)	,
(	45365	)	,
(	45351	)	,
(	45337	)	,
(	45323	)	,
(	45310	)	,
(	45296	)	,
(	45282	)	,
(	45268	)	,
(	45254	)	,
(	45241	)	,
(	45227	)	,
(	45213	)	,
(	45199	)	,
(	45186	)	,
(	45172	)	,
(	45158	)	,
(	45144	)	,
(	45130	)	,
(	45117	)	,
(	45103	)	,
(	45089	)	,
(	45075	)	,
(	45061	)	,
(	45048	)	,
(	45034	)	,
(	45020	)	,
(	45006	)	,
(	44992	)	,
(	44979	)	,
(	44965	)	,
(	44951	)	,
(	44937	)	,
(	44924	)	,
(	44910	)	,
(	44896	)	,
(	44882	)	,
(	44868	)	,
(	44855	)	,
(	44841	)	,
(	44827	)	,
(	44813	)	,
(	44799	)	,
(	44786	)	,
(	44772	)	,
(	44758	)	,
(	44744	)	,
(	44730	)	,
(	44717	)	,
(	44703	)	,
(	44689	)	,
(	44675	)	,
(	44662	)	,
(	44648	)	,
(	44634	)	,
(	44620	)	,
(	44606	)	,
(	44593	)	,
(	44579	)	,
(	44565	)	,
(	44551	)	,
(	44537	)	,
(	44524	)	,
(	44510	)	,
(	44496	)	,
(	44482	)	,
(	44469	)	,
(	44455	)	,
(	44441	)	,
(	44427	)	,
(	44413	)	,
(	44400	)	,
(	44386	)	,
(	44372	)	,
(	44358	)	,
(	44344	)	,
(	44331	)	,
(	44317	)	,
(	44303	)	,
(	44289	)	,
(	44275	)	,
(	44262	)	,
(	44248	)	,
(	44234	)	,
(	44220	)	,
(	44207	)	,
(	44193	)	,
(	44179	)	,
(	44165	)	,
(	44151	)	,
(	44138	)	,
(	44124	)	,
(	44110	)	,
(	44096	)	,
(	44082	)	,
(	44069	)	,
(	44055	)	,
(	44041	)	,
(	44027	)	,
(	44013	)	,
(	44000	)	,
(	43986	)	,
(	43972	)	,
(	43958	)	,
(	43945	)	,
(	43931	)	,
(	43917	)	,
(	43903	)	,
(	43889	)	,
(	43876	)	,
(	43862	)	,
(	43848	)	,
(	43834	)	,
(	43820	)	,
(	43807	)	,
(	43793	)	,
(	43779	)	,
(	43765	)	,
(	43751	)	,
(	43738	)	,
(	43724	)	,
(	43710	)	,
(	43696	)	,
(	43683	)	,
(	43669	)	,
(	43655	)	,
(	43641	)	,
(	43627	)	,
(	43614	)	,
(	43600	)	,
(	43586	)	,
(	43572	)	,
(	43558	)	,
(	43545	)	,
(	43531	)	,
(	43517	)	,
(	43503	)	,
(	43489	)	,
(	43476	)	,
(	43462	)	,
(	43448	)	,
(	43434	)	,
(	43421	)	,
(	43407	)	,
(	43393	)	,
(	43379	)	,
(	43365	)	,
(	43352	)	,
(	43338	)	,
(	43324	)	,
(	43310	)	,
(	43296	)	,
(	43283	)	,
(	43269	)	,
(	43255	)	,
(	43241	)	,
(	43227	)	,
(	43214	)	,
(	43200	)	,
(	43186	)	,
(	43172	)	,
(	43159	)	,
(	43145	)	,
(	43131	)	,
(	43117	)	,
(	43103	)	,
(	43090	)	,
(	43076	)	,
(	43062	)	,
(	43048	)	,
(	43034	)	,
(	43021	)	,
(	43007	)	,
(	42993	)	,
(	42979	)	,
(	42965	)	,
(	42952	)	,
(	42938	)	,
(	42924	)	,
(	42910	)	,
(	42897	)	,
(	42883	)	,
(	42869	)	,
(	42855	)	,
(	42841	)	,
(	42828	)	,
(	42814	)	,
(	42800	)	,
(	42786	)	,
(	42772	)	,
(	42759	)	,
(	42745	)	,
(	42731	)	,
(	42717	)	,
(	42704	)	,
(	42690	)	,
(	42676	)	,
(	42662	)	,
(	42648	)	,
(	42635	)	,
(	42621	)	,
(	42607	)	,
(	42593	)	,
(	42579	)	,
(	42566	)	,
(	42552	)	,
(	42538	)	,
(	42524	)	,
(	42510	)	,
(	42497	)	,
(	42483	)	,
(	42469	)	,
(	42455	)	,
(	42442	)	,
(	42428	)	,
(	42414	)	,
(	42400	)	,
(	42386	)	,
(	42373	)	,
(	42359	)	,
(	42345	)	,
(	42331	)	,
(	42317	)	,
(	42304	)	,
(	42290	)	,
(	42276	)	,
(	42262	)	,
(	42248	)	,
(	42235	)	,
(	42221	)	,
(	42207	)	,
(	42193	)	,
(	42180	)	,
(	42166	)	,
(	42152	)	,
(	42138	)	,
(	42124	)	,
(	42111	)	,
(	42097	)	,
(	42083	)	,
(	42069	)	,
(	42055	)	,
(	42042	)	,
(	42028	)	,
(	42014	)	,
(	42000	)	,
(	41986	)	,
(	41973	)	,
(	41959	)	,
(	41945	)	,
(	41931	)	,
(	41918	)	,
(	41904	)	,
(	41890	)	,
(	41876	)	,
(	41862	)	,
(	41849	)	,
(	41835	)	,
(	41821	)	,
(	41807	)	,
(	41793	)	,
(	41780	)	,
(	41766	)	,
(	41752	)	,
(	41738	)	,
(	41724	)	,
(	41711	)	,
(	41697	)	,
(	41683	)	,
(	41669	)	,
(	41656	)	,
(	41642	)	,
(	41628	)	,
(	41614	)	,
(	41600	)	,
(	41587	)	,
(	41573	)	,
(	41559	)	,
(	41545	)	,
(	41531	)	,
(	41518	)	,
(	41504	)	,
(	41490	)	,
(	41476	)	,
(	41462	)	,
(	41449	)	,
(	41435	)	,
(	41421	)	,
(	41407	)	,
(	41394	)	,
(	41380	)	,
(	41366	)	,
(	41352	)	,
(	41338	)	,
(	41325	)	,
(	41311	)	,
(	41297	)	,
(	41283	)	,
(	41269	)	,
(	41256	)	,
(	41242	)	,
(	41228	)	,
(	41214	)	,
(	41201	)	,
(	41187	)	,
(	41173	)	,
(	41159	)	,
(	41145	)	,
(	41132	)	,
(	41118	)	,
(	41104	)	,
(	41090	)	,
(	41076	)	,
(	41063	)	,
(	41049	)	,
(	41035	)	,
(	41021	)	,
(	41007	)	,
(	40994	)	,
(	40980	)	,
(	40966	)	,
(	40952	)	,
(	40939	)	,
(	40925	)	,
(	40911	)	,
(	40897	)	,
(	40883	)	,
(	40870	)	,
(	40856	)	,
(	40842	)	,
(	40828	)	,
(	40814	)	,
(	40801	)	,
(	40787	)	,
(	40773	)	,
(	40759	)	,
(	40745	)	,
(	40732	)	,
(	40718	)	,
(	40704	)	,
(	40690	)	,
(	40677	)	,
(	40663	)	,
(	40649	)	,
(	40635	)	,
(	40621	)	,
(	40608	)	,
(	40594	)	,
(	40580	)	,
(	40566	)	,
(	40552	)	,
(	40539	)	,
(	40525	)	,
(	40511	)	,
(	40497	)	,
(	40483	)	,
(	40470	)	,
(	40456	)	,
(	40442	)	,
(	40428	)	,
(	40415	)	,
(	40401	)	,
(	40387	)	,
(	40373	)	,
(	40359	)	,
(	40346	)	,
(	40332	)	,
(	40318	)	,
(	40304	)	,
(	40290	)	,
(	40277	)	,
(	40263	)	,
(	40249	)	,
(	40235	)	,
(	40221	)	,
(	40208	)	,
(	40194	)	,
(	40180	)	,
(	40166	)	,
(	40153	)	,
(	40139	)	,
(	40125	)	,
(	40111	)	,
(	40097	)	,
(	40084	)	,
(	40070	)	,
(	40056	)	,
(	40042	)	,
(	40028	)	,
(	40015	)	,
(	40001	)	,
(	39987	)	,
(	39973	)	,
(	39959	)	,
(	39946	)	,
(	39932	)	,
(	39918	)	,
(	39904	)	,
(	39891	)	,
(	39877	)	,
(	39863	)	,
(	39849	)	,
(	39835	)	,
(	39822	)	,
(	39808	)	,
(	39794	)	,
(	39780	)	,
(	39766	)	,
(	39753	)	,
(	39739	)	,
(	39725	)	,
(	39711	)	,
(	39698	)	,
(	39684	)	,
(	39670	)	,
(	39656	)	,
(	39642	)	,
(	39629	)	,
(	39615	)	,
(	39601	)	,
(	39587	)	,
(	39573	)	,
(	39560	)	,
(	39546	)	,
(	39532	)	,
(	39518	)	,
(	39504	)	,
(	39491	)	,
(	39477	)	,
(	39463	)	,
(	39449	)	,
(	39436	)	,
(	39422	)	,
(	39408	)	,
(	39394	)	,
(	39380	)	,
(	39367	)	,
(	39353	)	,
(	39339	)	,
(	39325	)	,
(	39311	)	,
(	39298	)	,
(	39284	)	,
(	39270	)	,
(	39256	)	,
(	39242	)	,
(	39229	)	,
(	39215	)	,
(	39201	)	,
(	39187	)	,
(	39174	)	,
(	39160	)	,
(	39146	)	,
(	39132	)	,
(	39118	)	,
(	39105	)	,
(	39091	)	,
(	39077	)	,
(	39063	)	,
(	39049	)	,
(	39036	)	,
(	39022	)	,
(	39008	)	,
(	38994	)	,
(	38980	)	,
(	38967	)	,
(	38953	)	,
(	38939	)	,
(	38925	)	,
(	38912	)	,
(	38898	)	,
(	38884	)	,
(	38870	)	,
(	38856	)	,
(	38843	)	,
(	38829	)	,
(	38815	)	,
(	38801	)	,
(	38787	)	,
(	38774	)	,
(	38760	)	,
(	38746	)	,
(	38732	)	,
(	38718	)	,
(	38705	)	,
(	38691	)	,
(	38677	)	,
(	38663	)	,
(	38650	)	,
(	38636	)	,
(	38622	)	,
(	38608	)	,
(	38594	)	,
(	38581	)	,
(	38567	)	,
(	38553	)	,
(	38539	)	,
(	38525	)	,
(	38512	)	,
(	38498	)	,
(	38484	)	,
(	38470	)	,
(	38456	)	,
(	38443	)	,
(	38429	)	,
(	38415	)	,
(	38401	)	,
(	38388	)	,
(	38374	)	,
(	38360	)	,
(	38346	)	,
(	38332	)	,
(	38319	)	,
(	38305	)	,
(	38291	)	,
(	38277	)	,
(	38263	)	,
(	38250	)	,
(	38236	)	,
(	38222	)	,
(	38208	)	,
(	38195	)	,
(	38181	)	,
(	38167	)	,
(	38153	)	,
(	38139	)	,
(	38126	)	,
(	38112	)	,
(	38098	)	,
(	38084	)	,
(	38070	)	,
(	38057	)	,
(	38043	)	,
(	38029	)	,
(	38015	)	,
(	38001	)	,
(	37988	)	,
(	37974	)	,
(	37960	)	,
(	37946	)	,
(	37933	)	,
(	37919	)	,
(	37905	)	,
(	37891	)	,
(	37877	)	,
(	37864	)	,
(	37850	)	,
(	37836	)	,
(	37822	)	,
(	37808	)	,
(	37795	)	,
(	37781	)	,
(	37767	)	,
(	37753	)	,
(	37739	)	,
(	37726	)	,
(	37712	)	,
(	37698	)	,
(	37684	)	,
(	37671	)	,
(	37657	)	,
(	37643	)	,
(	37629	)	,
(	37615	)	,
(	37602	)	,
(	37588	)	,
(	37574	)	,
(	37560	)	,
(	37546	)	,
(	37533	)	,
(	37519	)	,
(	37505	)	,
(	37491	)	,
(	37477	)	,
(	37464	)	,
(	37450	)	,
(	37436	)	,
(	37422	)	,
(	37409	)	,
(	37395	)	,
(	37381	)	,
(	37367	)	,
(	37353	)	,
(	37340	)	,
(	37326	)	,
(	37312	)	,
(	37298	)	,
(	37284	)	,
(	37271	)	,
(	37257	)	,
(	37243	)	,
(	37229	)	,
(	37215	)	,
(	37202	)	,
(	37188	)	,
(	37174	)	,
(	37160	)	,
(	37147	)	,
(	37133	)	,
(	37119	)	,
(	37105	)	,
(	37091	)	,
(	37078	)	,
(	37064	)	,
(	37050	)	,
(	37036	)	,
(	37022	)	,
(	37009	)	,
(	36995	)	,
(	36981	)	,
(	36967	)	,
(	36953	)	,
(	36940	)	,
(	36926	)	,
(	36912	)	,
(	36898	)	,
(	36885	)	,
(	36871	)	,
(	36857	)	,
(	36843	)	,
(	36829	)	,
(	36816	)	,
(	36802	)	,
(	36788	)	,
(	36774	)	,
(	36760	)	,
(	36747	)	,
(	36733	)	,
(	36719	)	,
(	36705	)	,
(	36692	)	,
(	36678	)	,
(	36664	)	,
(	36650	)	,
(	36636	)	,
(	36623	)	,
(	36609	)	,
(	36595	)	,
(	36581	)	,
(	36567	)	,
(	36554	)	,
(	36540	)	,
(	36526	)	,
(	36512	)	,
(	36498	)	,
(	36485	)	,
(	36471	)	,
(	36457	)	,
(	36443	)	,
(	36430	)	,
(	36416	)	,
(	36402	)	,
(	36388	)	,
(	36374	)	,
(	36361	)	,
(	36347	)	,
(	36333	)	,
(	36319	)	,
(	36305	)	,
(	36292	)	,
(	36278	)	,
(	36264	)	,
(	36250	)	,
(	36236	)	,
(	36223	)	,
(	36209	)	,
(	36195	)	,
(	36181	)	,
(	36168	)	,
(	36154	)	,
(	36140	)	,
(	36126	)	,
(	36112	)	,
(	36099	)	,
(	36085	)	,
(	36071	)	,
(	36057	)	,
(	36043	)	,
(	36030	)	,
(	36016	)	,
(	36002	)	,
(	35988	)	,
(	35974	)	,
(	35961	)	,
(	35947	)	,
(	35933	)	,
(	35919	)	,
(	35906	)	,
(	35892	)	,
(	35878	)	,
(	35864	)	,
(	35850	)	,
(	35837	)	,
(	35823	)	,
(	35809	)	,
(	35795	)	,
(	35781	)	,
(	35768	)	,
(	35754	)	,
(	35740	)	,
(	35726	)	,
(	35712	)	,
(	35699	)	,
(	35685	)	,
(	35671	)	,
(	35657	)	,
(	35644	)	,
(	35630	)	,
(	35616	)	,
(	35602	)	,
(	35588	)	,
(	35575	)	,
(	35561	)	,
(	35547	)	,
(	35533	)	,
(	35519	)	,
(	35506	)	,
(	35492	)	,
(	35478	)	,
(	35464	)	,
(	35450	)	,
(	35437	)	,
(	35423	)	,
(	35409	)	,
(	35395	)	,
(	35382	)	,
(	35368	)	,
(	35354	)	,
(	35340	)	,
(	35326	)	,
(	35313	)	,
(	35299	)	,
(	35285	)	,
(	35271	)	,
(	35257	)	,
(	35244	)	,
(	35230	)	,
(	35216	)	,
(	35202	)	,
(	35189	)	,
(	35175	)	,
(	35161	)	,
(	35147	)	,
(	35133	)	,
(	35120	)	,
(	35106	)	,
(	35092	)	,
(	35078	)	,
(	35064	)	,
(	35051	)	,
(	35037	)	,
(	35023	)	,
(	35009	)	,
(	34995	)	,
(	34982	)	,
(	34968	)	,
(	34954	)	,
(	34940	)	,
(	34927	)	,
(	34913	)	,
(	34899	)	,
(	34885	)	,
(	34871	)	,
(	34858	)	,
(	34844	)	,
(	34830	)	,
(	34816	)	,
(	34802	)	,
(	34789	)	,
(	34775	)	,
(	34761	)	,
(	34747	)	,
(	34733	)	,
(	34720	)	,
(	34706	)	,
(	34692	)	,
(	34678	)	,
(	34665	)	,
(	34651	)	,
(	34637	)	,
(	34623	)	,
(	34609	)	,
(	34596	)	,
(	34582	)	,
(	34568	)	,
(	34554	)	,
(	34540	)	,
(	34527	)	,
(	34513	)	,
(	34499	)	,
(	34485	)	,
(	34471	)	,
(	34458	)	,
(	34444	)	,
(	34430	)	,
(	34416	)	,
(	34403	)	,
(	34389	)	,
(	34375	)	,
(	34361	)	,
(	34347	)	,
(	34334	)	,
(	34320	)	,
(	34306	)	,
(	34292	)	,
(	34278	)	,
(	34265	)	,
(	34251	)	,
(	34237	)	,
(	34223	)	,
(	34209	)	,
(	34196	)	,
(	34182	)	,
(	34168	)	,
(	34154	)	,
(	34141	)	,
(	34127	)	,
(	34113	)	,
(	34099	)	,
(	34085	)	,
(	34072	)	,
(	34058	)	,
(	34044	)	,
(	34030	)	,
(	34016	)	,
(	34003	)	,
(	33989	)	,
(	33975	)	,
(	33961	)	,
(	33947	)	,
(	33934	)	,
(	33920	)	,
(	33906	)	,
(	33892	)	,
(	33879	)	,
(	33865	)	,
(	33851	)	,
(	33837	)	,
(	33823	)	,
(	33810	)	,
(	33796	)	,
(	33782	)	,
(	33768	)	,
(	33754	)	,
(	33741	)	,
(	33727	)	,
(	33713	)	,
(	33699	)	,
(	33686	)	,
(	33672	)	,
(	33658	)	,
(	33644	)	,
(	33630	)	,
(	33617	)	,
(	33603	)	,
(	33589	)	,
(	33575	)	,
(	33561	)	,
(	33548	)	,
(	33534	)	,
(	33520	)	,
(	33506	)	,
(	33492	)	,
(	33479	)	,
(	33465	)	,
(	33451	)	,
(	33437	)	,
(	33424	)	,
(	33410	)	,
(	33396	)	,
(	33382	)	,
(	33368	)	,
(	33355	)	,
(	33341	)	,
(	33327	)	,
(	33313	)	,
(	33299	)	,
(	33286	)	,
(	33272	)	,
(	33258	)	,
(	33244	)	,
(	33230	)	,
(	33217	)	,
(	33203	)	,
(	33189	)	,
(	33175	)	,
(	33162	)	,
(	33148	)	,
(	33134	)	,
(	33120	)	,
(	33106	)	,
(	33093	)	,
(	33079	)	,
(	33065	)	,
(	33051	)	,
(	33037	)	,
(	33024	)	,
(	33010	)	,
(	32996	)	,
(	32982	)	,
(	32968	)	,
(	32955	)	,
(	32941	)	,
(	32927	)	,
(	32913	)	,
(	32900	)	,
(	32886	)	,
(	32872	)	,
(	32858	)	,
(	32844	)	,
(	32831	)	,
(	32817	)	,
(	32803	)	,
(	32789	)	,
(	32775	)	,
(	32762	)	,
(	32748	)	,
(	32734	)	,
(	32720	)	,
(	32706	)	,
(	32693	)	,
(	32679	)	,
(	32665	)	,
(	32651	)	,
(	32638	)	,
(	32624	)	,
(	32610	)	,
(	32596	)	,
(	32582	)	,
(	32569	)	,
(	32555	)	,
(	32541	)	,
(	32527	)	,
(	32513	)	,
(	32500	)	,
(	32486	)	,
(	32472	)	,
(	32458	)	,
(	32444	)	,
(	32431	)	,
(	32417	)	,
(	32403	)	,
(	32389	)	,
(	32376	)	,
(	32362	)	,
(	32348	)	,
(	32334	)	,
(	32320	)	,
(	32307	)	,
(	32293	)	,
(	32279	)	,
(	32265	)	,
(	32251	)	,
(	32238	)	,
(	32224	)	,
(	32210	)	,
(	32196	)	,
(	32183	)	,
(	32169	)	,
(	32155	)	,
(	32141	)	,
(	32127	)	,
(	32114	)	,
(	32100	)	,
(	32086	)	,
(	32072	)	,
(	32058	)	,
(	32045	)	,
(	32031	)	,
(	32017	)	,
(	32003	)	,
(	31989	)	,
(	31976	)	,
(	31962	)	,
(	31948	)	,
(	31934	)	,
(	31921	)	,
(	31907	)	,
(	31893	)	,
(	31879	)	,
(	31865	)	,
(	31852	)	,
(	31838	)	,
(	31824	)	,
(	31810	)	,
(	31796	)	,
(	31783	)	,
(	31769	)	,
(	31755	)	,
(	31741	)	,
(	31727	)	,
(	31714	)	,
(	31700	)	,
(	31686	)	,
(	31672	)	,
(	31659	)	,
(	31645	)	,
(	31631	)	,
(	31617	)	,
(	31603	)	,
(	31590	)	,
(	31576	)	,
(	31562	)	,
(	31548	)	,
(	31534	)	,
(	31521	)	,
(	31507	)	,
(	31493	)	,
(	31479	)	,
(	31465	)	,
(	31452	)	,
(	31438	)	,
(	31424	)	,
(	31410	)	,
(	31397	)	,
(	31383	)	,
(	31369	)	,
(	31355	)	,
(	31341	)	,
(	31328	)	,
(	31314	)	,
(	31300	)	,
(	31286	)	,
(	31272	)	,
(	31259	)	,
(	31245	)	,
(	31231	)	,
(	31217	)	,
(	31203	)	,
(	31190	)	,
(	31176	)	,
(	31162	)	,
(	31148	)	,
(	31135	)	,
(	31121	)	,
(	31107	)	,
(	31093	)	,
(	31079	)	,
(	31066	)	,
(	31052	)	,
(	31038	)	,
(	31024	)	,
(	31010	)	,
(	30997	)	,
(	30983	)	,
(	30969	)	,
(	30955	)	,
(	30941	)	,
(	30928	)	,
(	30914	)	,
(	30900	)	,
(	30886	)	,
(	30873	)	,
(	30859	)	,
(	30845	)	,
(	30831	)	,
(	30817	)	,
(	30804	)	,
(	30790	)	,
(	30776	)	,
(	30762	)	,
(	30748	)	,
(	30735	)	,
(	30721	)	,
(	30707	)	,
(	30693	)	,
(	30680	)	,
(	30666	)	,
(	30652	)	,
(	30638	)	,
(	30624	)	,
(	30611	)	,
(	30597	)	,
(	30583	)	,
(	30569	)	,
(	30555	)	,
(	30542	)	,
(	30528	)	,
(	30514	)	,
(	30500	)	,
(	30486	)	,
(	30473	)	,
(	30459	)	,
(	30445	)	,
(	30431	)	,
(	30418	)	,
(	30404	)	,
(	30390	)	,
(	30376	)	,
(	30362	)	,
(	30349	)	,
(	30335	)	,
(	30321	)	,
(	30307	)	,
(	30293	)	,
(	30280	)	,
(	30266	)	,
(	30252	)	,
(	30238	)	,
(	30224	)	,
(	30211	)	,
(	30197	)	,
(	30183	)	,
(	30169	)	,
(	30156	)	,
(	30142	)	,
(	30128	)	,
(	30114	)	,
(	30100	)	,
(	30087	)	,
(	30073	)	,
(	30059	)	,
(	30045	)	,
(	30031	)	,
(	30018	)	,
(	30004	)	,
(	29990	)	,
(	29976	)	,
(	29962	)	,
(	29949	)	,
(	29935	)	,
(	29921	)	,
(	29907	)	,
(	29894	)	,
(	29880	)	,
(	29866	)	,
(	29852	)	,
(	29838	)	,
(	29825	)	,
(	29811	)	,
(	29797	)	,
(	29783	)	,
(	29769	)	,
(	29756	)	,
(	29742	)	,
(	29728	)	,
(	29714	)	,
(	29700	)	,
(	29687	)	,
(	29673	)	,
(	29659	)	,
(	29645	)	,
(	29632	)	,
(	29618	)	,
(	29604	)	,
(	29590	)	,
(	29576	)	,
(	29563	)	,
(	29549	)	,
(	29535	)	,
(	29521	)	,
(	29507	)	,
(	29494	)	,
(	29480	)	,
(	29466	)	,
(	29452	)	,
(	29438	)	,
(	29425	)	,
(	29411	)	,
(	29397	)	,
(	29383	)	,
(	29370	)	,
(	29356	)	,
(	29342	)	,
(	29328	)	,
(	29314	)	,
(	29301	)	,
(	29287	)	,
(	29273	)	,
(	29259	)	,
(	29245	)	,
(	29232	)	,
(	29218	)	,
(	29204	)	,
(	29190	)	,
(	29176	)	,
(	29163	)	,
(	29149	)	,
(	29135	)	,
(	29121	)	,
(	29108	)	,
(	29094	)	,
(	29080	)	,
(	29066	)	,
(	29052	)	,
(	29039	)	,
(	29025	)	,
(	29011	)	,
(	28997	)	,
(	28983	)	,
(	28970	)	,
(	28956	)	,
(	28942	)	,
(	28928	)	,
(	28915	)	,
(	28901	)	,
(	28887	)	,
(	28873	)	,
(	28859	)	,
(	28846	)	,
(	28832	)	,
(	28818	)	,
(	28804	)	,
(	28790	)	,
(	28777	)	,
(	28763	)	,
(	28749	)	,
(	28735	)	,
(	28721	)	,
(	28708	)	,
(	28694	)	,
(	28680	)	,
(	28666	)	,
(	28653	)	,
(	28639	)	,
(	28625	)	,
(	28611	)	,
(	28597	)	,
(	28584	)	,
(	28570	)	,
(	28556	)	,
(	28542	)	,
(	28528	)	,
(	28515	)	,
(	28501	)	,
(	28487	)	,
(	28473	)	,
(	28459	)	,
(	28446	)	,
(	28432	)	,
(	28418	)	,
(	28404	)	,
(	28391	)	,
(	28377	)	,
(	28363	)	,
(	28349	)	,
(	28335	)	,
(	28322	)	,
(	28308	)	,
(	28294	)	,
(	28280	)	,
(	28266	)	,
(	28253	)	,
(	28239	)	,
(	28225	)	,
(	28211	)	,
(	28197	)	,
(	28184	)	,
(	28170	)	,
(	28156	)	,
(	28142	)	,
(	28129	)	,
(	28115	)	,
(	28101	)	,
(	28087	)	,
(	28073	)	,
(	28060	)	,
(	28046	)	,
(	28032	)	,
(	28018	)	,
(	28004	)	,
(	27991	)	,
(	27977	)	,
(	27963	)	,
(	27949	)	,
(	27935	)	,
(	27922	)	,
(	27908	)	,
(	27894	)	,
(	27880	)	,
(	27867	)	,
(	27853	)	,
(	27839	)	,
(	27825	)	,
(	27811	)	,
(	27798	)	,
(	27784	)	,
(	27770	)	,
(	27756	)	,
(	27742	)	,
(	27729	)	,
(	27715	)	,
(	27701	)	,
(	27687	)	,
(	27673	)	,
(	27660	)	,
(	27646	)	,
(	27632	)	,
(	27618	)	,
(	27605	)	,
(	27591	)	,
(	27577	)	,
(	27563	)	,
(	27549	)	,
(	27536	)	,
(	27522	)	,
(	27508	)	,
(	27494	)	,
(	27480	)	,
(	27467	)	,
(	27453	)	,
(	27439	)	,
(	27425	)	,
(	27412	)	,
(	27398	)	,
(	27384	)	,
(	27370	)	,
(	27356	)	,
(	27343	)	,
(	27329	)	,
(	27315	)	,
(	27301	)	,
(	27287	)	,
(	27274	)	,
(	27260	)	,
(	27246	)	,
(	27232	)	,
(	27218	)	,
(	27205	)	,
(	27191	)	,
(	27177	)	,
(	27163	)	,
(	27150	)	,
(	27136	)	,
(	27122	)	,
(	27108	)	,
(	27094	)	,
(	27081	)	,
(	27067	)	,
(	27053	)	,
(	27039	)	,
(	27025	)	,
(	27012	)	,
(	26998	)	,
(	26984	)	,
(	26970	)	,
(	26956	)	,
(	26943	)	,
(	26929	)	,
(	26915	)	,
(	26901	)	,
(	26888	)	,
(	26874	)	,
(	26860	)	,
(	26846	)	,
(	26832	)	,
(	26819	)	,
(	26805	)	,
(	26791	)	,
(	26777	)	,
(	26763	)	,
(	26750	)	,
(	26736	)	,
(	26722	)	,
(	26708	)	,
(	26694	)	,
(	26681	)	,
(	26667	)	,
(	26653	)	,
(	26639	)	,
(	26626	)	,
(	26612	)	,
(	26598	)	,
(	26584	)	,
(	26570	)	,
(	26557	)	,
(	26543	)	,
(	26529	)	,
(	26515	)	,
(	26501	)	,
(	26488	)	,
(	26474	)	,
(	26460	)	,
(	26446	)	,
(	26432	)	,
(	26419	)	,
(	26405	)	,
(	26391	)	,
(	26377	)	,
(	26364	)	,
(	26350	)	,
(	26336	)	,
(	26322	)	,
(	26308	)	,
(	26295	)	,
(	26281	)	,
(	26267	)	,
(	26253	)	,
(	26239	)	,
(	26226	)	,
(	26212	)	,
(	26198	)	,
(	26184	)	,
(	26170	)	,
(	26157	)	,
(	26143	)	,
(	26129	)	,
(	26115	)	,
(	26102	)	,
(	26088	)	,
(	26074	)	,
(	26060	)	,
(	26046	)	,
(	26033	)	,
(	26019	)	,
(	26005	)	,
(	25991	)	,
(	25977	)	,
(	25964	)	,
(	25950	)	,
(	25936	)	,
(	25922	)	,
(	25909	)	,
(	25895	)	,
(	25881	)	,
(	25867	)	,
(	25853	)	,
(	25840	)	,
(	25826	)	,
(	25812	)	,
(	25798	)	,
(	25784	)	,
(	25771	)	,
(	25757	)	,
(	25743	)	,
(	25729	)	,
(	25715	)	,
(	25702	)	,
(	25688	)	,
(	25674	)	,
(	25660	)	,
(	25647	)	,
(	25633	)	,
(	25619	)	,
(	25605	)	,
(	25591	)	,
(	25578	)	,
(	25564	)	,
(	25550	)	,
(	25536	)	,
(	25522	)	,
(	25509	)	,
(	25495	)	,
(	25481	)	,
(	25467	)	,
(	25453	)	,
(	25440	)	,
(	25426	)	,
(	25412	)	,
(	25398	)	,
(	25385	)	,
(	25371	)	,
(	25357	)	,
(	25343	)	,
(	25329	)	,
(	25316	)	,
(	25302	)	,
(	25288	)	,
(	25274	)	,
(	25260	)	,
(	25247	)	,
(	25233	)	,
(	25219	)	,
(	25205	)	,
(	25191	)	,
(	25178	)	,
(	25164	)	,
(	25150	)	,
(	25136	)	,
(	25123	)	,
(	25109	)	,
(	25095	)	,
(	25081	)	,
(	25067	)	,
(	25054	)	,
(	25040	)	,
(	25026	)	,
(	25012	)	,
(	24998	)	,
(	24985	)	,
(	24971	)	,
(	24957	)	,
(	24943	)	,
(	24929	)	,
(	24916	)	,
(	24902	)	,
(	24888	)	,
(	24874	)	,
(	24861	)	,
(	24847	)	,
(	24833	)	,
(	24819	)	,
(	24805	)	,
(	24792	)	,
(	24778	)	,
(	24764	)	,
(	24750	)	,
(	24736	)	,
(	24723	)	,
(	24709	)	,
(	24695	)	,
(	24681	)	,
(	24667	)	,
(	24654	)	,
(	24640	)	,
(	24626	)	,
(	24612	)	,
(	24599	)	,
(	24585	)	,
(	24571	)	,
(	24557	)	,
(	24543	)	,
(	24530	)	,
(	24516	)	,
(	24502	)	,
(	24488	)	,
(	24474	)	,
(	24461	)	,
(	24447	)	,
(	24433	)	,
(	24419	)	,
(	24406	)	,
(	24392	)	,
(	24378	)	,
(	24364	)	,
(	24350	)	,
(	24337	)	,
(	24323	)	,
(	24309	)	,
(	24295	)	,
(	24281	)	,
(	24268	)	,
(	24254	)	,
(	24240	)	,
(	24226	)	,
(	24212	)	,
(	24199	)	,
(	24185	)	,
(	24171	)	,
(	24157	)	,
(	24144	)	,
(	24130	)	,
(	24116	)	,
(	24102	)	,
(	24088	)	,
(	24075	)	,
(	24061	)	,
(	24047	)	,
(	24033	)	,
(	24019	)	,
(	24006	)	,
(	23992	)	,
(	23978	)	,
(	23964	)	,
(	23950	)	,
(	23937	)	,
(	23923	)	,
(	23909	)	,
(	23895	)	,
(	23882	)	,
(	23868	)	,
(	23854	)	,
(	23840	)	,
(	23826	)	,
(	23813	)	,
(	23799	)	,
(	23785	)	,
(	23771	)	,
(	23757	)	,
(	23744	)	,
(	23730	)	,
(	23716	)	,
(	23702	)	,
(	23688	)	,
(	23675	)	,
(	23661	)	,
(	23647	)	,
(	23633	)	,
(	23620	)	,
(	23606	)	,
(	23592	)	,
(	23578	)	,
(	23564	)	,
(	23551	)	,
(	23537	)	,
(	23523	)	,
(	23509	)	,
(	23495	)	,
(	23482	)	,
(	23468	)	,
(	23454	)	,
(	23440	)	,
(	23426	)	,
(	23413	)	,
(	23399	)	,
(	23385	)	,
(	23371	)	,
(	23358	)	,
(	23344	)	,
(	23330	)	,
(	23316	)	,
(	23302	)	,
(	23289	)	,
(	23275	)	,
(	23261	)	,
(	23247	)	,
(	23233	)	,
(	23220	)	,
(	23206	)	,
(	23192	)	,
(	23178	)	,
(	23164	)	,
(	23151	)	,
(	23137	)	,
(	23123	)	,
(	23109	)	,
(	23096	)	,
(	23082	)	,
(	23068	)	,
(	23054	)	,
(	23040	)	,
(	23027	)	,
(	23013	)	,
(	22999	)	,
(	22985	)	,
(	22971	)	,
(	22958	)	,
(	22944	)	,
(	22930	)	,
(	22916	)	,
(	22903	)	,
(	22889	)	,
(	22875	)	,
(	22861	)	,
(	22847	)	,
(	22834	)	,
(	22820	)	,
(	22806	)	,
(	22792	)	,
(	22778	)	,
(	22765	)	,
(	22751	)	,
(	22737	)	,
(	22723	)	,
(	22709	)	,
(	22696	)	,
(	22682	)	,
(	22668	)	,
(	22654	)	,
(	22641	)	,
(	22627	)	,
(	22613	)	,
(	22599	)	,
(	22585	)	,
(	22572	)	,
(	22558	)	,
(	22544	)	,
(	22530	)	,
(	22516	)	,
(	22503	)	,
(	22489	)	,
(	22475	)	,
(	22461	)	,
(	22447	)	,
(	22434	)	,
(	22420	)	,
(	22406	)	,
(	22392	)	,
(	22379	)	,
(	22365	)	,
(	22351	)	,
(	22337	)	,
(	22323	)	,
(	22310	)	,
(	22296	)	,
(	22282	)	,
(	22268	)	,
(	22254	)	,
(	22241	)	,
(	22227	)	,
(	22213	)	,
(	22199	)	,
(	22185	)	,
(	22172	)	,
(	22158	)	,
(	22144	)	,
(	22130	)	,
(	22117	)	,
(	22103	)	,
(	22089	)	,
(	22075	)	,
(	22061	)	,
(	22048	)	,
(	22034	)	,
(	22020	)	,
(	22006	)	,
(	21992	)	,
(	21979	)	,
(	21965	)	,
(	21951	)	,
(	21937	)	,
(	21923	)	,
(	21910	)	,
(	21896	)	,
(	21882	)	,
(	21868	)	,
(	21855	)	,
(	21841	)	,
(	21827	)	,
(	21813	)	,
(	21799	)	,
(	21786	)	,
(	21772	)	,
(	21758	)	,
(	21744	)	,
(	21730	)	,
(	21717	)	,
(	21703	)	,
(	21689	)	,
(	21675	)	,
(	21661	)	,
(	21648	)	,
(	21634	)	,
(	21620	)	,
(	21606	)	,
(	21593	)	,
(	21579	)	,
(	21565	)	,
(	21551	)	,
(	21537	)	,
(	21524	)	,
(	21510	)	,
(	21496	)	,
(	21482	)	,
(	21468	)	,
(	21455	)	,
(	21441	)	,
(	21427	)	,
(	21413	)	,
(	21400	)	,
(	21386	)	,
(	21372	)	,
(	21358	)	,
(	21344	)	,
(	21331	)	,
(	21317	)	,
(	21303	)	,
(	21289	)	,
(	21275	)	,
(	21262	)	,
(	21248	)	,
(	21234	)	,
(	21220	)	,
(	21206	)	,
(	21193	)	,
(	21179	)	,
(	21165	)	,
(	21151	)	,
(	21138	)	,
(	21124	)	,
(	21110	)	,
(	21096	)	,
(	21082	)	,
(	21069	)	,
(	21055	)	,
(	21041	)	,
(	21027	)	,
(	21013	)	,
(	21000	)	,
(	20986	)	,
(	20972	)	,
(	20958	)	,
(	20944	)	,
(	20931	)	,
(	20917	)	,
(	20903	)	,
(	20889	)	,
(	20876	)	,
(	20862	)	,
(	20848	)	,
(	20834	)	,
(	20820	)	,
(	20807	)	,
(	20793	)	,
(	20779	)	,
(	20765	)	,
(	20751	)	,
(	20738	)	,
(	20724	)	,
(	20710	)	,
(	20696	)	,
(	20682	)	,
(	20669	)	,
(	20655	)	,
(	20641	)	,
(	20627	)	,
(	20614	)	,
(	20600	)	,
(	20586	)	,
(	20572	)	,
(	20558	)	,
(	20545	)	,
(	20531	)	,
(	20517	)	,
(	20503	)	,
(	20489	)	,
(	20476	)	,
(	20462	)	,
(	20448	)	,
(	20434	)	,
(	20420	)	,
(	20407	)	,
(	20393	)	,
(	20379	)	,
(	20365	)	,
(	20352	)	,
(	20338	)	,
(	20324	)	,
(	20310	)	,
(	20296	)	,
(	20283	)	,
(	20269	)	,
(	20255	)	,
(	20241	)	,
(	20227	)	,
(	20214	)	,
(	20200	)	,
(	20186	)	,
(	20172	)	,
(	20158	)	,
(	20145	)	,
(	20131	)	,
(	20117	)	,
(	20103	)	,
(	20090	)	,
(	20076	)	,
(	20062	)	,
(	20048	)	,
(	20034	)	,
(	20021	)	,
(	20007	)	,
(	19993	)	,
(	19979	)	,
(	19965	)	,
(	19952	)	,
(	19938	)	,
(	19924	)	,
(	19910	)	,
(	19897	)	,
(	19883	)	,
(	19869	)	,
(	19855	)	,
(	19841	)	,
(	19828	)	,
(	19814	)	,
(	19800	)	,
(	19786	)	,
(	19772	)	,
(	19759	)	,
(	19745	)	,
(	19731	)	,
(	19717	)	,
(	19703	)	,
(	19690	)	,
(	19676	)	,
(	19662	)	,
(	19648	)	,
(	19635	)	,
(	19621	)	,
(	19607	)	,
(	19593	)	,
(	19579	)	,
(	19566	)	,
(	19552	)	,
(	19538	)	,
(	19524	)	,
(	19510	)	,
(	19497	)	,
(	19483	)	,
(	19469	)	,
(	19455	)	,
(	19441	)	,
(	19428	)	,
(	19414	)	,
(	19400	)	,
(	19386	)	,
(	19373	)	,
(	19359	)	,
(	19345	)	,
(	19331	)	,
(	19317	)	,
(	19304	)	,
(	19290	)	,
(	19276	)	,
(	19262	)	,
(	19248	)	,
(	19235	)	,
(	19221	)	,
(	19207	)	,
(	19193	)	,
(	19179	)	,
(	19166	)	,
(	19152	)	,
(	19138	)	,
(	19124	)	,
(	19111	)	,
(	19097	)	,
(	19083	)	,
(	19069	)	,
(	19055	)	,
(	19042	)	,
(	19028	)	,
(	19014	)	,
(	19000	)	,
(	18986	)	,
(	18973	)	,
(	18959	)	,
(	18945	)	,
(	18931	)	,
(	18917	)	,
(	18904	)	,
(	18890	)	,
(	18876	)	,
(	18862	)	,
(	18849	)	,
(	18835	)	,
(	18821	)	,
(	18807	)	,
(	18793	)	,
(	18780	)	,
(	18766	)	,
(	18752	)	,
(	18738	)	,
(	18724	)	,
(	18711	)	,
(	18697	)	,
(	18683	)	,
(	18669	)	,
(	18655	)	,
(	18642	)	,
(	18628	)	,
(	18614	)	,
(	18600	)	,
(	18587	)	,
(	18573	)	,
(	18559	)	,
(	18545	)	,
(	18531	)	,
(	18518	)	,
(	18504	)	,
(	18490	)	,
(	18476	)	,
(	18462	)	,
(	18449	)	,
(	18435	)	,
(	18421	)	,
(	18407	)	,
(	18394	)	,
(	18380	)	,
(	18366	)	,
(	18352	)	,
(	18338	)	,
(	18325	)	,
(	18311	)	,
(	18297	)	,
(	18283	)	,
(	18269	)	,
(	18256	)	,
(	18242	)	,
(	18228	)	,
(	18214	)	,
(	18200	)	,
(	18187	)	,
(	18173	)	,
(	18159	)	,
(	18145	)	,
(	18132	)	,
(	18118	)	,
(	18104	)	,
(	18090	)	,
(	18076	)	,
(	18063	)	,
(	18049	)	,
(	18035	)	,
(	18021	)	,
(	18007	)	,
(	17994	)	,
(	17980	)	,
(	17966	)	,
(	17952	)	,
(	17938	)	,
(	17925	)	,
(	17911	)	,
(	17897	)	,
(	17883	)	,
(	17870	)	,
(	17856	)	,
(	17842	)	,
(	17828	)	,
(	17814	)	,
(	17801	)	,
(	17787	)	,
(	17773	)	,
(	17759	)	,
(	17745	)	,
(	17732	)	,
(	17718	)	,
(	17704	)	,
(	17690	)	,
(	17676	)	,
(	17663	)	,
(	17649	)	,
(	17635	)	,
(	17621	)	,
(	17608	)	,
(	17594	)	,
(	17580	)	,
(	17566	)	,
(	17552	)	,
(	17539	)	,
(	17525	)	,
(	17511	)	,
(	17497	)	,
(	17483	)	,
(	17470	)	,
(	17456	)	,
(	17442	)	,
(	17428	)	,
(	17414	)	,
(	17401	)	,
(	17387	)	,
(	17373	)	,
(	17359	)	,
(	17346	)	,
(	17332	)	,
(	17318	)	,
(	17304	)	,
(	17290	)	,
(	17277	)	,
(	17263	)	,
(	17249	)	,
(	17235	)	,
(	17221	)	,
(	17208	)	,
(	17194	)	,
(	17180	)	,
(	17166	)	,
(	17152	)	,
(	17139	)	,
(	17125	)	,
(	17111	)	,
(	17097	)	,
(	17084	)	,
(	17070	)	,
(	17056	)	,
(	17042	)	,
(	17028	)	,
(	17015	)	,
(	17001	)	,
(	16987	)	,
(	16973	)	,
(	16959	)	,
(	16946	)	,
(	16932	)	,
(	16918	)	,
(	16904	)	,
(	16891	)	,
(	16877	)	,
(	16863	)	,
(	16849	)	,
(	16835	)	,
(	16822	)	,
(	16808	)	,
(	16794	)	,
(	16780	)	,
(	16766	)	,
(	16753	)	,
(	16739	)	,
(	16725	)	,
(	16711	)	,
(	16697	)	,
(	16684	)	,
(	16670	)	,
(	16656	)	,
(	16642	)	,
(	16629	)	,
(	16615	)	,
(	16601	)	,
(	16587	)	,
(	16573	)	,
(	16560	)	,
(	16546	)	,
(	16532	)	,
(	16518	)	,
(	16504	)	,
(	16491	)	,
(	16477	)	,
(	16463	)	,
(	16449	)	,
(	16435	)	,
(	16422	)	,
(	16408	)	,
(	16394	)	,
(	16380	)	,
(	16367	)	,
(	16353	)	,
(	16339	)	,
(	16325	)	,
(	16311	)	,
(	16298	)	,
(	16284	)	,
(	16270	)	,
(	16256	)	,
(	16242	)	,
(	16229	)	,
(	16215	)	,
(	16201	)	,
(	16187	)	,
(	16173	)	,
(	16160	)	,
(	16146	)	,
(	16132	)	,
(	16118	)	,
(	16105	)	,
(	16091	)	,
(	16077	)	,
(	16063	)	,
(	16049	)	,
(	16036	)	,
(	16022	)	,
(	16008	)	,
(	15994	)	,
(	15980	)	,
(	15967	)	,
(	15953	)	,
(	15939	)	,
(	15925	)	,
(	15911	)	,
(	15898	)	,
(	15884	)	,
(	15870	)	,
(	15856	)	,
(	15843	)	,
(	15829	)	,
(	15815	)	,
(	15801	)	,
(	15787	)	,
(	15774	)	,
(	15760	)	,
(	15746	)	,
(	15732	)	,
(	15718	)	,
(	15705	)	,
(	15691	)	,
(	15677	)	,
(	15663	)	,
(	15649	)	,
(	15636	)	,
(	15622	)	,
(	15608	)	,
(	15594	)	,
(	15581	)	,
(	15567	)	,
(	15553	)	,
(	15539	)	,
(	15525	)	,
(	15512	)	,
(	15498	)	,
(	15484	)	,
(	15470	)	,
(	15456	)	,
(	15443	)	,
(	15429	)	,
(	15415	)	,
(	15401	)	,
(	15387	)	,
(	15374	)	,
(	15360	)	,
(	15346	)	,
(	15332	)	,
(	15319	)	,
(	15305	)	,
(	15291	)	,
(	15277	)	,
(	15263	)	,
(	15250	)	,
(	15236	)	,
(	15222	)	,
(	15208	)	,
(	15194	)	,
(	15181	)	,
(	15167	)	,
(	15153	)	,
(	15139	)	,
(	15126	)	,
(	15112	)	,
(	15098	)	,
(	15084	)	,
(	15070	)	,
(	15057	)	,
(	15043	)	,
(	15029	)	,
(	15015	)	,
(	15001	)	,
(	14988	)	,
(	14974	)	,
(	14960	)	,
(	14946	)	,
(	14932	)	,
(	14919	)	,
(	14905	)	,
(	14891	)	,
(	14877	)	,
(	14864	)	,
(	14850	)	,
(	14836	)	,
(	14822	)	,
(	14808	)	,
(	14795	)	,
(	14781	)	,
(	14767	)	,
(	14753	)	,
(	14739	)	,
(	14726	)	,
(	14712	)	,
(	14698	)	,
(	14684	)	,
(	14670	)	,
(	14657	)	,
(	14643	)	,
(	14629	)	,
(	14615	)	,
(	14602	)	,
(	14588	)	,
(	14574	)	,
(	14560	)	,
(	14546	)	,
(	14533	)	,
(	14519	)	,
(	14505	)	,
(	14491	)	,
(	14477	)	,
(	14464	)	,
(	14450	)	,
(	14436	)	,
(	14422	)	,
(	14408	)	,
(	14395	)	,
(	14381	)	,
(	14367	)	,
(	14353	)	,
(	14340	)	,
(	14326	)	,
(	14312	)	,
(	14298	)	,
(	14284	)	,
(	14271	)	,
(	14257	)	,
(	14243	)	,
(	14229	)	,
(	14215	)	,
(	14202	)	,
(	14188	)	,
(	14174	)	,
(	14160	)	,
(	14146	)	,
(	14133	)	,
(	14119	)	,
(	14105	)	,
(	14091	)	,
(	14078	)	,
(	14064	)	,
(	14050	)	,
(	14036	)	,
(	14022	)	,
(	14009	)	,
(	13995	)	,
(	13981	)	,
(	13967	)	,
(	13953	)	,
(	13940	)	,
(	13926	)	,
(	13912	)	,
(	13898	)	,
(	13884	)	,
(	13871	)	,
(	13857	)	,
(	13843	)	,
(	13829	)	,
(	13816	)	,
(	13802	)	,
(	13788	)	,
(	13774	)	,
(	13760	)	,
(	13747	)	,
(	13733	)	,
(	13719	)	,
(	13705	)	,
(	13691	)	,
(	13678	)	,
(	13664	)	,
(	13650	)	,
(	13636	)	,
(	13623	)	,
(	13609	)	,
(	13595	)	,
(	13581	)	,
(	13567	)	,
(	13554	)	,
(	13540	)	,
(	13526	)	,
(	13512	)	,
(	13498	)	,
(	13485	)	,
(	13471	)	,
(	13457	)	,
(	13443	)	,
(	13429	)	,
(	13416	)	,
(	13402	)	,
(	13388	)	,
(	13374	)	,
(	13361	)	,
(	13347	)	,
(	13333	)	,
(	13319	)	,
(	13305	)	,
(	13292	)	,
(	13278	)	,
(	13264	)	,
(	13250	)	,
(	13236	)	,
(	13223	)	,
(	13209	)	,
(	13195	)	,
(	13181	)	,
(	13167	)	,
(	13154	)	,
(	13140	)	,
(	13126	)	,
(	13112	)	,
(	13099	)	,
(	13085	)	,
(	13071	)	,
(	13057	)	,
(	13043	)	,
(	13030	)	,
(	13016	)	,
(	13002	)	,
(	12988	)	,
(	12974	)	,
(	12961	)	,
(	12947	)	,
(	12933	)	,
(	12919	)	,
(	12905	)	,
(	12892	)	,
(	12878	)	,
(	12864	)	,
(	12850	)	,
(	12837	)	,
(	12823	)	,
(	12809	)	,
(	12795	)	,
(	12781	)	,
(	12768	)	,
(	12754	)	,
(	12740	)	,
(	12726	)	,
(	12712	)	,
(	12699	)	,
(	12685	)	,
(	12671	)	,
(	12657	)	,
(	12643	)	,
(	12630	)	,
(	12616	)	,
(	12602	)	,
(	12588	)	,
(	12575	)	,
(	12561	)	,
(	12547	)	,
(	12533	)	,
(	12519	)	,
(	12506	)	,
(	12492	)	,
(	12478	)	,
(	12464	)	,
(	12450	)	,
(	12437	)	,
(	12423	)	,
(	12409	)	,
(	12395	)	,
(	12381	)	,
(	12368	)	,
(	12354	)	,
(	12340	)	,
(	12326	)	,
(	12313	)	,
(	12299	)	,
(	12285	)	,
(	12271	)	,
(	12257	)	,
(	12244	)	,
(	12230	)	,
(	12216	)	,
(	12202	)	,
(	12188	)	,
(	12175	)	,
(	12161	)	,
(	12147	)	,
(	12133	)	,
(	12120	)	,
(	12106	)	,
(	12092	)	,
(	12078	)	,
(	12064	)	,
(	12051	)	,
(	12037	)	,
(	12023	)	,
(	12009	)	,
(	11995	)	,
(	11982	)	,
(	11968	)	,
(	11954	)	,
(	11940	)	,
(	11926	)	,
(	11913	)	,
(	11899	)	,
(	11885	)	,
(	11871	)	,
(	11858	)	,
(	11844	)	,
(	11830	)	,
(	11816	)	,
(	11802	)	,
(	11789	)	,
(	11775	)	,
(	11761	)	,
(	11747	)	,
(	11733	)	,
(	11720	)	,
(	11706	)	,
(	11692	)	,
(	11678	)	,
(	11664	)	,
(	11651	)	,
(	11637	)	,
(	11623	)	,
(	11609	)	,
(	11596	)	,
(	11582	)	,
(	11568	)	,
(	11554	)	,
(	11540	)	,
(	11527	)	,
(	11513	)	,
(	11499	)	,
(	11485	)	,
(	11471	)	,
(	11458	)	,
(	11444	)	,
(	11430	)	,
(	11416	)	,
(	11402	)	,
(	11389	)	,
(	11375	)	,
(	11361	)	,
(	11347	)	,
(	11334	)	,
(	11320	)	,
(	11306	)	,
(	11292	)	,
(	11278	)	,
(	11265	)	,
(	11251	)	,
(	11237	)	,
(	11223	)	,
(	11209	)	,
(	11196	)	,
(	11182	)	,
(	11168	)	,
(	11154	)	,
(	11140	)	,
(	11127	)	,
(	11113	)	,
(	11099	)	,
(	11085	)	,
(	11072	)	,
(	11058	)	,
(	11044	)	,
(	11030	)	,
(	11016	)	,
(	11003	)	,
(	10989	)	,
(	10975	)	,
(	10961	)	,
(	10947	)	,
(	10934	)	,
(	10920	)	,
(	10906	)	,
(	10892	)	,
(	10878	)	,
(	10865	)	,
(	10851	)	,
(	10837	)	,
(	10823	)	,
(	10810	)	,
(	10796	)	,
(	10782	)	,
(	10768	)	,
(	10754	)	,
(	10741	)	,
(	10727	)	,
(	10713	)	,
(	10699	)	,
(	10685	)	,
(	10672	)	,
(	10658	)	,
(	10644	)	,
(	10630	)	,
(	10617	)	,
(	10603	)	,
(	10589	)	,
(	10575	)	,
(	10561	)	,
(	10548	)	,
(	10534	)	,
(	10520	)	,
(	10506	)	,
(	10492	)	,
(	10479	)	,
(	10465	)	,
(	10451	)	,
(	10437	)	,
(	10423	)	,
(	10410	)	,
(	10396	)	,
(	10382	)	,
(	10368	)	,
(	10355	)	,
(	10341	)	,
(	10327	)	,
(	10313	)	,
(	10299	)	,
(	10286	)	,
(	10272	)	,
(	10258	)	,
(	10244	)	,
(	10230	)	,
(	10217	)	,
(	10203	)	,
(	10189	)	,
(	10175	)	,
(	10161	)	,
(	10148	)	,
(	10134	)	,
(	10120	)	,
(	10106	)	,
(	10093	)	,
(	10079	)	,
(	10065	)	,
(	10051	)	,
(	10037	)	,
(	10024	)	,
(	10010	)	,
(	9996	)	,
(	9982	)	,
(	9968	)	,
(	9955	)	,
(	9941	)	,
(	9927	)	,
(	9913	)	,
(	9899	)	,
(	9886	)	,
(	9872	)	,
(	9858	)	,
(	9844	)	,
(	9831	)	,
(	9817	)	,
(	9803	)	,
(	9789	)	,
(	9775	)	,
(	9762	)	,
(	9748	)	,
(	9734	)	,
(	9720	)	,
(	9706	)	,
(	9693	)	,
(	9679	)	,
(	9665	)	,
(	9651	)	,
(	9637	)	,
(	9624	)	,
(	9610	)	,
(	9596	)	,
(	9582	)	,
(	9569	)	,
(	9555	)	,
(	9541	)	,
(	9527	)	,
(	9513	)	,
(	9500	)	,
(	9486	)	,
(	9472	)	,
(	9458	)	,
(	9444	)	,
(	9431	)	,
(	9417	)	,
(	9403	)	,
(	9389	)	,
(	9375	)	,
(	9362	)	,
(	9348	)	,
(	9334	)	,
(	9320	)	,
(	9307	)	,
(	9293	)	,
(	9279	)	,
(	9265	)	,
(	9251	)	,
(	9238	)	,
(	9224	)	,
(	9210	)	,
(	9196	)	,
(	9182	)	,
(	9169	)	,
(	9155	)	,
(	9141	)	,
(	9127	)	,
(	9114	)	,
(	9100	)	,
(	9086	)	,
(	9072	)	,
(	9058	)	,
(	9045	)	,
(	9031	)	,
(	9017	)	,
(	9003	)	,
(	8989	)	,
(	8976	)	,
(	8962	)	,
(	8948	)	,
(	8934	)	,
(	8920	)	,
(	8907	)	,
(	8893	)	,
(	8879	)	,
(	8865	)	,
(	8852	)	,
(	8838	)	,
(	8824	)	,
(	8810	)	,
(	8796	)	,
(	8783	)	,
(	8769	)	,
(	8755	)	,
(	8741	)	,
(	8727	)	,
(	8714	)	,
(	8700	)	,
(	8686	)	

);

end package LUT_flashing_pkg;