library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_flashing_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 5414) of integer;
constant d2freq_LUT : array_1d := (

(	-7903	)	,
(	-7867	)	,
(	-7830	)	,
(	-7794	)	,
(	-7757	)	,
(	-7721	)	,
(	-7684	)	,
(	-7648	)	,
(	-7612	)	,
(	-7575	)	,
(	-7539	)	,
(	-7502	)	,
(	-7466	)	,
(	-7429	)	,
(	-7393	)	,
(	-7356	)	,
(	-7320	)	,
(	-7284	)	,
(	-7247	)	,
(	-7211	)	,
(	-7174	)	,
(	-7138	)	,
(	-7101	)	,
(	-7065	)	,
(	-7028	)	,
(	-6992	)	,
(	-6955	)	,
(	-6919	)	,
(	-6883	)	,
(	-6846	)	,
(	-6810	)	,
(	-6773	)	,
(	-6737	)	,
(	-6700	)	,
(	-6664	)	,
(	-6627	)	,
(	-6591	)	,
(	-6554	)	,
(	-6518	)	,
(	-6482	)	,
(	-6445	)	,
(	-6409	)	,
(	-6372	)	,
(	-6336	)	,
(	-6299	)	,
(	-6263	)	,
(	-6226	)	,
(	-6190	)	,
(	-6154	)	,
(	-6117	)	,
(	-6081	)	,
(	-6044	)	,
(	-6008	)	,
(	-5971	)	,
(	-5935	)	,
(	-5898	)	,
(	-5862	)	,
(	-5825	)	,
(	-5789	)	,
(	-5753	)	,
(	-5716	)	,
(	-5680	)	,
(	-5643	)	,
(	-5607	)	,
(	-5570	)	,
(	-5534	)	,
(	-5497	)	,
(	-5461	)	,
(	-5424	)	,
(	-5388	)	,
(	-5352	)	,
(	-5315	)	,
(	-5279	)	,
(	-5242	)	,
(	-5206	)	,
(	-5169	)	,
(	-5133	)	,
(	-5096	)	,
(	-5060	)	,
(	-5023	)	,
(	-4987	)	,
(	-4951	)	,
(	-4914	)	,
(	-4878	)	,
(	-4841	)	,
(	-4805	)	,
(	-4768	)	,
(	-4732	)	,
(	-4695	)	,
(	-4659	)	,
(	-4623	)	,
(	-4586	)	,
(	-4550	)	,
(	-4513	)	,
(	-4477	)	,
(	-4440	)	,
(	-4404	)	,
(	-4367	)	,
(	-4331	)	,
(	-4294	)	,
(	-4258	)	,
(	-4222	)	,
(	-4185	)	,
(	-4149	)	,
(	-4112	)	,
(	-4076	)	,
(	-4039	)	,
(	-4003	)	,
(	-3966	)	,
(	-3930	)	,
(	-3893	)	,
(	-3857	)	,
(	-3821	)	,
(	-3784	)	,
(	-3748	)	,
(	-3711	)	,
(	-3675	)	,
(	-3638	)	,
(	-3602	)	,
(	-3565	)	,
(	-3529	)	,
(	-3493	)	,
(	-3456	)	,
(	-3420	)	,
(	-3383	)	,
(	-3347	)	,
(	-3310	)	,
(	-3274	)	,
(	-3237	)	,
(	-3201	)	,
(	-3164	)	,
(	-3128	)	,
(	-3092	)	,
(	-3055	)	,
(	-3019	)	,
(	-2982	)	,
(	-2946	)	,
(	-2909	)	,
(	-2873	)	,
(	-2836	)	,
(	-2800	)	,
(	-2763	)	,
(	-2727	)	,
(	-2691	)	,
(	-2654	)	,
(	-2618	)	,
(	-2581	)	,
(	-2545	)	,
(	-2508	)	,
(	-2472	)	,
(	-2435	)	,
(	-2399	)	,
(	-2362	)	,
(	-2326	)	,
(	-2290	)	,
(	-2253	)	,
(	-2217	)	,
(	-2180	)	,
(	-2144	)	,
(	-2107	)	,
(	-2071	)	,
(	-2034	)	,
(	-1998	)	,
(	-1962	)	,
(	-1925	)	,
(	-1889	)	,
(	-1852	)	,
(	-1816	)	,
(	-1779	)	,
(	-1743	)	,
(	-1706	)	,
(	-1670	)	,
(	-1633	)	,
(	-1597	)	,
(	-1561	)	,
(	-1524	)	,
(	-1488	)	,
(	-1451	)	,
(	-1415	)	,
(	-1378	)	,
(	-1342	)	,
(	-1305	)	,
(	-1269	)	,
(	-1232	)	,
(	-1196	)	,
(	-1160	)	,
(	-1123	)	,
(	-1087	)	,
(	-1050	)	,
(	-1014	)	,
(	-977	)	,
(	-941	)	,
(	-904	)	,
(	-868	)	,
(	-832	)	,
(	-795	)	,
(	-759	)	,
(	-722	)	,
(	-686	)	,
(	-649	)	,
(	-613	)	,
(	-576	)	,
(	-540	)	,
(	-503	)	,
(	-467	)	,
(	-431	)	,
(	-394	)	,
(	-358	)	,
(	-321	)	,
(	-285	)	,
(	-248	)	,
(	-212	)	,
(	-175	)	,
(	-139	)	,
(	-102	)	,
(	-66	)	,
(	-30	)	,
(	7	)	,
(	43	)	,
(	80	)	,
(	116	)	,
(	153	)	,
(	189	)	,
(	226	)	,
(	262	)	,
(	298	)	,
(	335	)	,
(	371	)	,
(	408	)	,
(	444	)	,
(	481	)	,
(	517	)	,
(	554	)	,
(	590	)	,
(	627	)	,
(	663	)	,
(	699	)	,
(	736	)	,
(	772	)	,
(	809	)	,
(	845	)	,
(	882	)	,
(	918	)	,
(	955	)	,
(	991	)	,
(	1028	)	,
(	1064	)	,
(	1100	)	,
(	1137	)	,
(	1173	)	,
(	1210	)	,
(	1246	)	,
(	1283	)	,
(	1319	)	,
(	1356	)	,
(	1392	)	,
(	1429	)	,
(	1465	)	,
(	1501	)	,
(	1538	)	,
(	1574	)	,
(	1611	)	,
(	1647	)	,
(	1684	)	,
(	1720	)	,
(	1757	)	,
(	1793	)	,
(	1829	)	,
(	1866	)	,
(	1902	)	,
(	1939	)	,
(	1975	)	,
(	2012	)	,
(	2048	)	,
(	2085	)	,
(	2121	)	,
(	2158	)	,
(	2194	)	,
(	2230	)	,
(	2267	)	,
(	2303	)	,
(	2340	)	,
(	2376	)	,
(	2413	)	,
(	2449	)	,
(	2486	)	,
(	2522	)	,
(	2559	)	,
(	2595	)	,
(	2631	)	,
(	2668	)	,
(	2704	)	,
(	2741	)	,
(	2777	)	,
(	2814	)	,
(	2850	)	,
(	2887	)	,
(	2923	)	,
(	2959	)	,
(	2996	)	,
(	3032	)	,
(	3069	)	,
(	3105	)	,
(	3142	)	,
(	3178	)	,
(	3215	)	,
(	3251	)	,
(	3288	)	,
(	3324	)	,
(	3360	)	,
(	3397	)	,
(	3433	)	,
(	3470	)	,
(	3506	)	,
(	3543	)	,
(	3579	)	,
(	3616	)	,
(	3652	)	,
(	3689	)	,
(	3725	)	,
(	3761	)	,
(	3798	)	,
(	3834	)	,
(	3871	)	,
(	3907	)	,
(	3944	)	,
(	3980	)	,
(	4017	)	,
(	4053	)	,
(	4090	)	,
(	4126	)	,
(	4162	)	,
(	4199	)	,
(	4235	)	,
(	4272	)	,
(	4308	)	,
(	4345	)	,
(	4381	)	,
(	4418	)	,
(	4454	)	,
(	4490	)	,
(	4527	)	,
(	4563	)	,
(	4600	)	,
(	4636	)	,
(	4673	)	,
(	4709	)	,
(	4746	)	,
(	4782	)	,
(	4819	)	,
(	4855	)	,
(	4891	)	,
(	4928	)	,
(	4964	)	,
(	5001	)	,
(	5037	)	,
(	5074	)	,
(	5110	)	,
(	5147	)	,
(	5183	)	,
(	5220	)	,
(	5256	)	,
(	5292	)	,
(	5329	)	,
(	5365	)	,
(	5402	)	,
(	5438	)	,
(	5475	)	,
(	5511	)	,
(	5548	)	,
(	5584	)	,
(	5620	)	,
(	5657	)	,
(	5693	)	,
(	5730	)	,
(	5766	)	,
(	5803	)	,
(	5839	)	,
(	5876	)	,
(	5912	)	,
(	5949	)	,
(	5985	)	,
(	6021	)	,
(	6058	)	,
(	6094	)	,
(	6131	)	,
(	6167	)	,
(	6204	)	,
(	6240	)	,
(	6277	)	,
(	6313	)	,
(	6350	)	,
(	6386	)	,
(	6422	)	,
(	6459	)	,
(	6495	)	,
(	6532	)	,
(	6568	)	,
(	6605	)	,
(	6641	)	,
(	6678	)	,
(	6714	)	,
(	6751	)	,
(	6787	)	,
(	6823	)	,
(	6860	)	,
(	6896	)	,
(	6933	)	,
(	6969	)	,
(	7006	)	,
(	7042	)	,
(	7079	)	,
(	7115	)	,
(	7151	)	,
(	7188	)	,
(	7224	)	,
(	7261	)	,
(	7297	)	,
(	7334	)	,
(	7370	)	,
(	7407	)	,
(	7443	)	,
(	7480	)	,
(	7516	)	,
(	7552	)	,
(	7589	)	,
(	7625	)	,
(	7662	)	,
(	7698	)	,
(	7735	)	,
(	7771	)	,
(	7808	)	,
(	7844	)	,
(	7881	)	,
(	7917	)	,
(	7953	)	,
(	7990	)	,
(	8026	)	,	  -- min distance = min period  = max frequnecy 
(	8063	)	,
(	8099	)	,
(	8136	)	,
(	8172	)	,
(	8209	)	,
(	8245	)	,
(	8281	)	,
(	8318	)	,
(	8354	)	,
(	8391	)	,
(	8427	)	,
(	8464	)	,
(	8500	)	,
(	8537	)	,
(	8573	)	,
(	8610	)	,
(	8646	)	,
(	8682	)	,
(	8719	)	,
(	8755	)	,
(	8792	)	,
(	8828	)	,
(	8865	)	,
(	8901	)	,
(	8938	)	,
(	8974	)	,
(	9011	)	,
(	9047	)	,
(	9083	)	,
(	9120	)	,
(	9156	)	,
(	9193	)	,
(	9229	)	,
(	9266	)	,
(	9302	)	,
(	9339	)	,
(	9375	)	,
(	9412	)	,
(	9448	)	,
(	9484	)	,
(	9521	)	,
(	9557	)	,
(	9594	)	,
(	9630	)	,
(	9667	)	,
(	9703	)	,
(	9740	)	,
(	9776	)	,
(	9812	)	,
(	9849	)	,
(	9885	)	,
(	9922	)	,
(	9958	)	,
(	9995	)	,
(	10031	)	,
(	10068	)	,
(	10104	)	,
(	10141	)	,
(	10177	)	,
(	10213	)	,
(	10250	)	,
(	10286	)	,
(	10323	)	,
(	10359	)	,
(	10396	)	,
(	10432	)	,
(	10469	)	,
(	10505	)	,
(	10542	)	,
(	10578	)	,
(	10614	)	,
(	10651	)	,
(	10687	)	,
(	10724	)	,
(	10760	)	,
(	10797	)	,
(	10833	)	,
(	10870	)	,
(	10906	)	,
(	10942	)	,
(	10979	)	,
(	11015	)	,
(	11052	)	,
(	11088	)	,
(	11125	)	,
(	11161	)	,
(	11198	)	,
(	11234	)	,
(	11271	)	,
(	11307	)	,
(	11343	)	,
(	11380	)	,
(	11416	)	,
(	11453	)	,
(	11489	)	,
(	11526	)	,
(	11562	)	,
(	11599	)	,
(	11635	)	,
(	11672	)	,
(	11708	)	,
(	11744	)	,
(	11781	)	,
(	11817	)	,
(	11854	)	,
(	11890	)	,
(	11927	)	,
(	11963	)	,
(	12000	)	,
(	12036	)	,
(	12072	)	,
(	12109	)	,
(	12145	)	,
(	12182	)	,
(	12218	)	,
(	12255	)	,
(	12291	)	,
(	12328	)	,
(	12364	)	,
(	12401	)	,
(	12437	)	,
(	12473	)	,
(	12510	)	,
(	12546	)	,
(	12583	)	,
(	12619	)	,
(	12656	)	,
(	12692	)	,
(	12729	)	,
(	12765	)	,
(	12802	)	,
(	12838	)	,
(	12874	)	,
(	12911	)	,
(	12947	)	,
(	12984	)	,
(	13020	)	,
(	13057	)	,
(	13093	)	,
(	13130	)	,
(	13166	)	,
(	13203	)	,
(	13239	)	,
(	13275	)	,
(	13312	)	,
(	13348	)	,
(	13385	)	,
(	13421	)	,
(	13458	)	,
(	13494	)	,
(	13531	)	,
(	13567	)	,
(	13603	)	,
(	13640	)	,
(	13676	)	,
(	13713	)	,
(	13749	)	,
(	13786	)	,
(	13822	)	,
(	13859	)	,
(	13895	)	,
(	13932	)	,
(	13968	)	,
(	14004	)	,
(	14041	)	,
(	14077	)	,
(	14114	)	,
(	14150	)	,
(	14187	)	,
(	14223	)	,
(	14260	)	,
(	14296	)	,
(	14333	)	,
(	14369	)	,
(	14405	)	,
(	14442	)	,
(	14478	)	,
(	14515	)	,
(	14551	)	,
(	14588	)	,
(	14624	)	,
(	14661	)	,
(	14697	)	,
(	14733	)	,
(	14770	)	,
(	14806	)	,
(	14843	)	,
(	14879	)	,
(	14916	)	,
(	14952	)	,
(	14989	)	,
(	15025	)	,
(	15062	)	,
(	15098	)	,
(	15134	)	,
(	15171	)	,
(	15207	)	,
(	15244	)	,
(	15280	)	,
(	15317	)	,
(	15353	)	,
(	15390	)	,
(	15426	)	,
(	15463	)	,
(	15499	)	,
(	15535	)	,
(	15572	)	,
(	15608	)	,
(	15645	)	,
(	15681	)	,
(	15718	)	,
(	15754	)	,
(	15791	)	,
(	15827	)	,
(	15864	)	,
(	15900	)	,
(	15936	)	,
(	15973	)	,
(	16009	)	,
(	16046	)	,
(	16082	)	,
(	16119	)	,
(	16155	)	,
(	16192	)	,
(	16228	)	,
(	16264	)	,
(	16301	)	,
(	16337	)	,
(	16374	)	,
(	16410	)	,
(	16447	)	,
(	16483	)	,
(	16520	)	,
(	16556	)	,
(	16593	)	,
(	16629	)	,
(	16665	)	,
(	16702	)	,
(	16738	)	,
(	16775	)	,
(	16811	)	,
(	16848	)	,
(	16884	)	,
(	16921	)	,
(	16957	)	,
(	16994	)	,
(	17030	)	,
(	17066	)	,
(	17103	)	,
(	17139	)	,
(	17176	)	,
(	17212	)	,
(	17249	)	,
(	17285	)	,
(	17322	)	,
(	17358	)	,
(	17394	)	,
(	17431	)	,
(	17467	)	,
(	17504	)	,
(	17540	)	,
(	17577	)	,
(	17613	)	,
(	17650	)	,
(	17686	)	,
(	17723	)	,
(	17759	)	,
(	17795	)	,
(	17832	)	,
(	17868	)	,
(	17905	)	,
(	17941	)	,
(	17978	)	,
(	18014	)	,
(	18051	)	,
(	18087	)	,
(	18124	)	,
(	18160	)	,
(	18196	)	,
(	18233	)	,
(	18269	)	,
(	18306	)	,
(	18342	)	,
(	18379	)	,
(	18415	)	,
(	18452	)	,
(	18488	)	,
(	18525	)	,
(	18561	)	,
(	18597	)	,
(	18634	)	,
(	18670	)	,
(	18707	)	,
(	18743	)	,
(	18780	)	,
(	18816	)	,
(	18853	)	,
(	18889	)	,
(	18925	)	,
(	18962	)	,
(	18998	)	,
(	19035	)	,
(	19071	)	,
(	19108	)	,
(	19144	)	,
(	19181	)	,
(	19217	)	,
(	19254	)	,
(	19290	)	,
(	19326	)	,
(	19363	)	,
(	19399	)	,
(	19436	)	,
(	19472	)	,
(	19509	)	,
(	19545	)	,
(	19582	)	,
(	19618	)	,
(	19655	)	,
(	19691	)	,
(	19727	)	,
(	19764	)	,
(	19800	)	,
(	19837	)	,
(	19873	)	,
(	19910	)	,
(	19946	)	,
(	19983	)	,
(	20019	)	,
(	20055	)	,
(	20092	)	,
(	20128	)	,
(	20165	)	,
(	20201	)	,
(	20238	)	,
(	20274	)	,
(	20311	)	,
(	20347	)	,
(	20384	)	,
(	20420	)	,
(	20456	)	,
(	20493	)	,
(	20529	)	,
(	20566	)	,
(	20602	)	,
(	20639	)	,
(	20675	)	,
(	20712	)	,
(	20748	)	,
(	20785	)	,
(	20821	)	,
(	20857	)	,
(	20894	)	,
(	20930	)	,
(	20967	)	,
(	21003	)	,
(	21040	)	,
(	21076	)	,
(	21113	)	,
(	21149	)	,
(	21185	)	,
(	21222	)	,
(	21258	)	,
(	21295	)	,
(	21331	)	,
(	21368	)	,
(	21404	)	,
(	21441	)	,
(	21477	)	,
(	21514	)	,
(	21550	)	,
(	21586	)	,
(	21623	)	,
(	21659	)	,
(	21696	)	,
(	21732	)	,
(	21769	)	,
(	21805	)	,
(	21842	)	,
(	21878	)	,
(	21915	)	,
(	21951	)	,
(	21987	)	,
(	22024	)	,
(	22060	)	,
(	22097	)	,
(	22133	)	,
(	22170	)	,
(	22206	)	,
(	22243	)	,
(	22279	)	,
(	22316	)	,
(	22352	)	,
(	22388	)	,
(	22425	)	,
(	22461	)	,
(	22498	)	,
(	22534	)	,
(	22571	)	,
(	22607	)	,
(	22644	)	,
(	22680	)	,
(	22716	)	,
(	22753	)	,
(	22789	)	,
(	22826	)	,
(	22862	)	,
(	22899	)	,
(	22935	)	,
(	22972	)	,
(	23008	)	,
(	23045	)	,
(	23081	)	,
(	23117	)	,
(	23154	)	,
(	23190	)	,
(	23227	)	,
(	23263	)	,
(	23300	)	,
(	23336	)	,
(	23373	)	,
(	23409	)	,
(	23446	)	,
(	23482	)	,
(	23518	)	,
(	23555	)	,
(	23591	)	,
(	23628	)	,
(	23664	)	,
(	23701	)	,
(	23737	)	,
(	23774	)	,
(	23810	)	,
(	23846	)	,
(	23883	)	,
(	23919	)	,
(	23956	)	,
(	23992	)	,
(	24029	)	,
(	24065	)	,
(	24102	)	,
(	24138	)	,
(	24175	)	,
(	24211	)	,
(	24247	)	,
(	24284	)	,
(	24320	)	,
(	24357	)	,
(	24393	)	,
(	24430	)	,
(	24466	)	,
(	24503	)	,
(	24539	)	,
(	24576	)	,
(	24612	)	,
(	24648	)	,
(	24685	)	,
(	24721	)	,
(	24758	)	,
(	24794	)	,
(	24831	)	,
(	24867	)	,
(	24904	)	,
(	24940	)	,
(	24977	)	,
(	25013	)	,
(	25049	)	,
(	25086	)	,
(	25122	)	,
(	25159	)	,
(	25195	)	,
(	25232	)	,
(	25268	)	,
(	25305	)	,
(	25341	)	,
(	25377	)	,
(	25414	)	,
(	25450	)	,
(	25487	)	,
(	25523	)	,
(	25560	)	,
(	25596	)	,
(	25633	)	,
(	25669	)	,
(	25706	)	,
(	25742	)	,
(	25778	)	,
(	25815	)	,
(	25851	)	,
(	25888	)	,
(	25924	)	,
(	25961	)	,
(	25997	)	,
(	26034	)	,
(	26070	)	,
(	26107	)	,
(	26143	)	,
(	26179	)	,
(	26216	)	,
(	26252	)	,
(	26289	)	,
(	26325	)	,
(	26362	)	,
(	26398	)	,
(	26435	)	,
(	26471	)	,
(	26507	)	,
(	26544	)	,
(	26580	)	,
(	26617	)	,
(	26653	)	,
(	26690	)	,
(	26726	)	,
(	26763	)	,
(	26799	)	,
(	26836	)	,
(	26872	)	,
(	26908	)	,
(	26945	)	,
(	26981	)	,
(	27018	)	,
(	27054	)	,
(	27091	)	,
(	27127	)	,
(	27164	)	,
(	27200	)	,
(	27237	)	,
(	27273	)	,
(	27309	)	,
(	27346	)	,
(	27382	)	,
(	27419	)	,
(	27455	)	,
(	27492	)	,
(	27528	)	,
(	27565	)	,
(	27601	)	,
(	27638	)	,
(	27674	)	,
(	27710	)	,
(	27747	)	,
(	27783	)	,
(	27820	)	,
(	27856	)	,
(	27893	)	,
(	27929	)	,
(	27966	)	,
(	28002	)	,
(	28038	)	,
(	28075	)	,
(	28111	)	,
(	28148	)	,
(	28184	)	,
(	28221	)	,
(	28257	)	,
(	28294	)	,
(	28330	)	,
(	28367	)	,
(	28403	)	,
(	28439	)	,
(	28476	)	,
(	28512	)	,
(	28549	)	,
(	28585	)	,
(	28622	)	,
(	28658	)	,
(	28695	)	,
(	28731	)	,
(	28768	)	,
(	28804	)	,
(	28840	)	,
(	28877	)	,
(	28913	)	,
(	28950	)	,
(	28986	)	,
(	29023	)	,
(	29059	)	,
(	29096	)	,
(	29132	)	,
(	29168	)	,
(	29205	)	,
(	29241	)	,
(	29278	)	,
(	29314	)	,
(	29351	)	,
(	29387	)	,
(	29424	)	,
(	29460	)	,
(	29497	)	,
(	29533	)	,
(	29569	)	,
(	29606	)	,
(	29642	)	,
(	29679	)	,
(	29715	)	,
(	29752	)	,
(	29788	)	,
(	29825	)	,
(	29861	)	,
(	29898	)	,
(	29934	)	,
(	29970	)	,
(	30007	)	,
(	30043	)	,
(	30080	)	,
(	30116	)	,
(	30153	)	,
(	30189	)	,
(	30226	)	,
(	30262	)	,
(	30298	)	,
(	30335	)	,
(	30371	)	,
(	30408	)	,
(	30444	)	,
(	30481	)	,
(	30517	)	,
(	30554	)	,
(	30590	)	,
(	30627	)	,
(	30663	)	,
(	30699	)	,
(	30736	)	,
(	30772	)	,
(	30809	)	,
(	30845	)	,
(	30882	)	,
(	30918	)	,
(	30955	)	,
(	30991	)	,
(	31028	)	,
(	31064	)	,
(	31100	)	,
(	31137	)	,
(	31173	)	,
(	31210	)	,
(	31246	)	,
(	31283	)	,
(	31319	)	,
(	31356	)	,
(	31392	)	,
(	31429	)	,
(	31465	)	,
(	31501	)	,
(	31538	)	,
(	31574	)	,
(	31611	)	,
(	31647	)	,
(	31684	)	,
(	31720	)	,
(	31757	)	,
(	31793	)	,
(	31829	)	,
(	31866	)	,
(	31902	)	,
(	31939	)	,
(	31975	)	,
(	32012	)	,
(	32048	)	,
(	32085	)	,
(	32121	)	,
(	32158	)	,
(	32194	)	,
(	32230	)	,
(	32267	)	,
(	32303	)	,
(	32340	)	,
(	32376	)	,
(	32413	)	,
(	32449	)	,
(	32486	)	,
(	32522	)	,
(	32559	)	,
(	32595	)	,
(	32631	)	,
(	32668	)	,
(	32704	)	,
(	32741	)	,
(	32777	)	,
(	32814	)	,
(	32850	)	,
(	32887	)	,
(	32923	)	,
(	32959	)	,
(	32996	)	,
(	33032	)	,
(	33069	)	,
(	33105	)	,
(	33142	)	,
(	33178	)	,
(	33215	)	,
(	33251	)	,
(	33288	)	,
(	33324	)	,
(	33360	)	,
(	33397	)	,
(	33433	)	,
(	33470	)	,
(	33506	)	,
(	33543	)	,
(	33579	)	,
(	33616	)	,
(	33652	)	,
(	33689	)	,
(	33725	)	,
(	33761	)	,
(	33798	)	,
(	33834	)	,
(	33871	)	,
(	33907	)	,
(	33944	)	,
(	33980	)	,
(	34017	)	,
(	34053	)	,
(	34090	)	,
(	34126	)	,
(	34162	)	,
(	34199	)	,
(	34235	)	,
(	34272	)	,
(	34308	)	,
(	34345	)	,
(	34381	)	,
(	34418	)	,
(	34454	)	,
(	34490	)	,
(	34527	)	,
(	34563	)	,
(	34600	)	,
(	34636	)	,
(	34673	)	,
(	34709	)	,
(	34746	)	,
(	34782	)	,
(	34819	)	,
(	34855	)	,
(	34891	)	,
(	34928	)	,
(	34964	)	,
(	35001	)	,
(	35037	)	,
(	35074	)	,
(	35110	)	,
(	35147	)	,
(	35183	)	,
(	35220	)	,
(	35256	)	,
(	35292	)	,
(	35329	)	,
(	35365	)	,
(	35402	)	,
(	35438	)	,
(	35475	)	,
(	35511	)	,
(	35548	)	,
(	35584	)	,
(	35620	)	,
(	35657	)	,
(	35693	)	,
(	35730	)	,
(	35766	)	,
(	35803	)	,
(	35839	)	,
(	35876	)	,
(	35912	)	,
(	35949	)	,
(	35985	)	,
(	36021	)	,
(	36058	)	,
(	36094	)	,
(	36131	)	,
(	36167	)	,
(	36204	)	,
(	36240	)	,
(	36277	)	,
(	36313	)	,
(	36350	)	,
(	36386	)	,
(	36422	)	,
(	36459	)	,
(	36495	)	,
(	36532	)	,
(	36568	)	,
(	36605	)	,
(	36641	)	,
(	36678	)	,
(	36714	)	,
(	36751	)	,
(	36787	)	,
(	36823	)	,
(	36860	)	,
(	36896	)	,
(	36933	)	,
(	36969	)	,
(	37006	)	,
(	37042	)	,
(	37079	)	,
(	37115	)	,
(	37151	)	,
(	37188	)	,
(	37224	)	,
(	37261	)	,
(	37297	)	,
(	37334	)	,
(	37370	)	,
(	37407	)	,
(	37443	)	,
(	37480	)	,
(	37516	)	,
(	37552	)	,
(	37589	)	,
(	37625	)	,
(	37662	)	,
(	37698	)	,
(	37735	)	,
(	37771	)	,
(	37808	)	,
(	37844	)	,
(	37881	)	,
(	37917	)	,
(	37953	)	,
(	37990	)	,
(	38026	)	,
(	38063	)	,
(	38099	)	,
(	38136	)	,
(	38172	)	,
(	38209	)	,
(	38245	)	,
(	38281	)	,
(	38318	)	,
(	38354	)	,
(	38391	)	,
(	38427	)	,
(	38464	)	,
(	38500	)	,
(	38537	)	,
(	38573	)	,
(	38610	)	,
(	38646	)	,
(	38682	)	,
(	38719	)	,
(	38755	)	,
(	38792	)	,
(	38828	)	,
(	38865	)	,
(	38901	)	,
(	38938	)	,
(	38974	)	,
(	39011	)	,
(	39047	)	,
(	39083	)	,
(	39120	)	,
(	39156	)	,
(	39193	)	,
(	39229	)	,
(	39266	)	,
(	39302	)	,
(	39339	)	,
(	39375	)	,
(	39411	)	,
(	39448	)	,
(	39484	)	,
(	39521	)	,
(	39557	)	,
(	39594	)	,
(	39630	)	,
(	39667	)	,
(	39703	)	,
(	39740	)	,
(	39776	)	,
(	39812	)	,
(	39849	)	,
(	39885	)	,
(	39922	)	,
(	39958	)	,
(	39995	)	,
(	40031	)	,
(	40068	)	,
(	40104	)	,
(	40141	)	,
(	40177	)	,
(	40213	)	,
(	40250	)	,
(	40286	)	,
(	40323	)	,
(	40359	)	,
(	40396	)	,
(	40432	)	,
(	40469	)	,
(	40505	)	,
(	40542	)	,
(	40578	)	,
(	40614	)	,
(	40651	)	,
(	40687	)	,
(	40724	)	,
(	40760	)	,
(	40797	)	,
(	40833	)	,
(	40870	)	,
(	40906	)	,
(	40942	)	,
(	40979	)	,
(	41015	)	,
(	41052	)	,
(	41088	)	,
(	41125	)	,
(	41161	)	,
(	41198	)	,
(	41234	)	,
(	41271	)	,
(	41307	)	,
(	41343	)	,
(	41380	)	,
(	41416	)	,
(	41453	)	,
(	41489	)	,
(	41526	)	,
(	41562	)	,
(	41599	)	,
(	41635	)	,
(	41672	)	,
(	41708	)	,
(	41744	)	,
(	41781	)	,
(	41817	)	,
(	41854	)	,
(	41890	)	,
(	41927	)	,
(	41963	)	,
(	42000	)	,
(	42036	)	,
(	42072	)	,
(	42109	)	,
(	42145	)	,
(	42182	)	,
(	42218	)	,
(	42255	)	,
(	42291	)	,
(	42328	)	,
(	42364	)	,
(	42401	)	,
(	42437	)	,
(	42473	)	,
(	42510	)	,
(	42546	)	,
(	42583	)	,
(	42619	)	,
(	42656	)	,
(	42692	)	,
(	42729	)	,
(	42765	)	,
(	42802	)	,
(	42838	)	,
(	42874	)	,
(	42911	)	,
(	42947	)	,
(	42984	)	,
(	43020	)	,
(	43057	)	,
(	43093	)	,
(	43130	)	,
(	43166	)	,
(	43203	)	,
(	43239	)	,
(	43275	)	,
(	43312	)	,
(	43348	)	,
(	43385	)	,
(	43421	)	,
(	43458	)	,
(	43494	)	,
(	43531	)	,
(	43567	)	,
(	43603	)	,
(	43640	)	,
(	43676	)	,
(	43713	)	,
(	43749	)	,
(	43786	)	,
(	43822	)	,
(	43859	)	,
(	43895	)	,
(	43932	)	,
(	43968	)	,
(	44004	)	,
(	44041	)	,
(	44077	)	,
(	44114	)	,
(	44150	)	,
(	44187	)	,
(	44223	)	,
(	44260	)	,
(	44296	)	,
(	44333	)	,
(	44369	)	,
(	44405	)	,
(	44442	)	,
(	44478	)	,
(	44515	)	,
(	44551	)	,
(	44588	)	,
(	44624	)	,
(	44661	)	,
(	44697	)	,
(	44733	)	,
(	44770	)	,
(	44806	)	,
(	44843	)	,
(	44879	)	,
(	44916	)	,
(	44952	)	,
(	44989	)	,
(	45025	)	,
(	45062	)	,
(	45098	)	,
(	45134	)	,
(	45171	)	,
(	45207	)	,
(	45244	)	,
(	45280	)	,
(	45317	)	,
(	45353	)	,
(	45390	)	,
(	45426	)	,
(	45463	)	,
(	45499	)	,
(	45535	)	,
(	45572	)	,
(	45608	)	,
(	45645	)	,
(	45681	)	,
(	45718	)	,
(	45754	)	,
(	45791	)	,
(	45827	)	,
(	45864	)	,
(	45900	)	,
(	45936	)	,
(	45973	)	,
(	46009	)	,
(	46046	)	,
(	46082	)	,
(	46119	)	,
(	46155	)	,
(	46192	)	,
(	46228	)	,
(	46264	)	,
(	46301	)	,
(	46337	)	,
(	46374	)	,
(	46410	)	,
(	46447	)	,
(	46483	)	,
(	46520	)	,
(	46556	)	,
(	46593	)	,
(	46629	)	,
(	46665	)	,
(	46702	)	,
(	46738	)	,
(	46775	)	,
(	46811	)	,
(	46848	)	,
(	46884	)	,
(	46921	)	,
(	46957	)	,
(	46994	)	,
(	47030	)	,
(	47066	)	,
(	47103	)	,
(	47139	)	,
(	47176	)	,
(	47212	)	,
(	47249	)	,
(	47285	)	,
(	47322	)	,
(	47358	)	,
(	47394	)	,
(	47431	)	,
(	47467	)	,
(	47504	)	,
(	47540	)	,
(	47577	)	,
(	47613	)	,
(	47650	)	,
(	47686	)	,
(	47723	)	,
(	47759	)	,
(	47795	)	,
(	47832	)	,
(	47868	)	,
(	47905	)	,
(	47941	)	,
(	47978	)	,
(	48014	)	,
(	48051	)	,
(	48087	)	,
(	48124	)	,
(	48160	)	,
(	48196	)	,
(	48233	)	,
(	48269	)	,
(	48306	)	,
(	48342	)	,
(	48379	)	,
(	48415	)	,
(	48452	)	,
(	48488	)	,
(	48524	)	,
(	48561	)	,
(	48597	)	,
(	48634	)	,
(	48670	)	,
(	48707	)	,
(	48743	)	,
(	48780	)	,
(	48816	)	,
(	48853	)	,
(	48889	)	,
(	48925	)	,
(	48962	)	,
(	48998	)	,
(	49035	)	,
(	49071	)	,
(	49108	)	,
(	49144	)	,
(	49181	)	,
(	49217	)	,
(	49254	)	,
(	49290	)	,
(	49326	)	,
(	49363	)	,
(	49399	)	,
(	49436	)	,
(	49472	)	,
(	49509	)	,
(	49545	)	,
(	49582	)	,
(	49618	)	,
(	49655	)	,
(	49691	)	,
(	49727	)	,
(	49764	)	,
(	49800	)	,
(	49837	)	,
(	49873	)	,
(	49910	)	,
(	49946	)	,
(	49983	)	,
(	50019	)	,
(	50055	)	,
(	50092	)	,
(	50128	)	,
(	50165	)	,
(	50201	)	,
(	50238	)	,
(	50274	)	,
(	50311	)	,
(	50347	)	,
(	50384	)	,
(	50420	)	,
(	50456	)	,
(	50493	)	,
(	50529	)	,
(	50566	)	,
(	50602	)	,
(	50639	)	,
(	50675	)	,
(	50712	)	,
(	50748	)	,
(	50785	)	,
(	50821	)	,
(	50857	)	,
(	50894	)	,
(	50930	)	,
(	50967	)	,
(	51003	)	,
(	51040	)	,
(	51076	)	,
(	51113	)	,
(	51149	)	,
(	51185	)	,
(	51222	)	,
(	51258	)	,
(	51295	)	,
(	51331	)	,
(	51368	)	,
(	51404	)	,
(	51441	)	,
(	51477	)	,
(	51514	)	,
(	51550	)	,
(	51586	)	,
(	51623	)	,
(	51659	)	,
(	51696	)	,
(	51732	)	,
(	51769	)	,
(	51805	)	,
(	51842	)	,
(	51878	)	,
(	51915	)	,
(	51951	)	,
(	51987	)	,
(	52024	)	,
(	52060	)	,
(	52097	)	,
(	52133	)	,
(	52170	)	,
(	52206	)	,
(	52243	)	,
(	52279	)	,
(	52316	)	,
(	52352	)	,
(	52388	)	,
(	52425	)	,
(	52461	)	,
(	52498	)	,
(	52534	)	,
(	52571	)	,
(	52607	)	,
(	52644	)	,
(	52680	)	,
(	52716	)	,
(	52753	)	,
(	52789	)	,
(	52826	)	,
(	52862	)	,
(	52899	)	,
(	52935	)	,
(	52972	)	,
(	53008	)	,
(	53045	)	,
(	53081	)	,
(	53117	)	,
(	53154	)	,
(	53190	)	,
(	53227	)	,
(	53263	)	,
(	53300	)	,
(	53336	)	,
(	53373	)	,
(	53409	)	,
(	53446	)	,
(	53482	)	,
(	53518	)	,
(	53555	)	,
(	53591	)	,
(	53628	)	,
(	53664	)	,
(	53701	)	,
(	53737	)	,
(	53774	)	,
(	53810	)	,
(	53846	)	,
(	53883	)	,
(	53919	)	,
(	53956	)	,
(	53992	)	,
(	54029	)	,
(	54065	)	,
(	54102	)	,
(	54138	)	,
(	54175	)	,
(	54211	)	,
(	54247	)	,
(	54284	)	,
(	54320	)	,
(	54357	)	,
(	54393	)	,
(	54430	)	,
(	54466	)	,
(	54503	)	,
(	54539	)	,
(	54576	)	,
(	54612	)	,
(	54648	)	,
(	54685	)	,
(	54721	)	,
(	54758	)	,
(	54794	)	,
(	54831	)	,
(	54867	)	,
(	54904	)	,
(	54940	)	,
(	54977	)	,
(	55013	)	,
(	55049	)	,
(	55086	)	,
(	55122	)	,
(	55159	)	,
(	55195	)	,
(	55232	)	,
(	55268	)	,
(	55305	)	,
(	55341	)	,
(	55377	)	,
(	55414	)	,
(	55450	)	,
(	55487	)	,
(	55523	)	,
(	55560	)	,
(	55596	)	,
(	55633	)	,
(	55669	)	,
(	55706	)	,
(	55742	)	,
(	55778	)	,
(	55815	)	,
(	55851	)	,
(	55888	)	,
(	55924	)	,
(	55961	)	,
(	55997	)	,
(	56034	)	,
(	56070	)	,
(	56107	)	,
(	56143	)	,
(	56179	)	,
(	56216	)	,
(	56252	)	,
(	56289	)	,
(	56325	)	,
(	56362	)	,
(	56398	)	,
(	56435	)	,
(	56471	)	,
(	56507	)	,
(	56544	)	,
(	56580	)	,
(	56617	)	,
(	56653	)	,
(	56690	)	,
(	56726	)	,
(	56763	)	,
(	56799	)	,
(	56836	)	,
(	56872	)	,
(	56908	)	,
(	56945	)	,
(	56981	)	,
(	57018	)	,
(	57054	)	,
(	57091	)	,
(	57127	)	,
(	57164	)	,
(	57200	)	,
(	57237	)	,
(	57273	)	,
(	57309	)	,
(	57346	)	,
(	57382	)	,
(	57419	)	,
(	57455	)	,
(	57492	)	,
(	57528	)	,
(	57565	)	,
(	57601	)	,
(	57637	)	,
(	57674	)	,
(	57710	)	,
(	57747	)	,
(	57783	)	,
(	57820	)	,
(	57856	)	,
(	57893	)	,
(	57929	)	,
(	57966	)	,
(	58002	)	,
(	58038	)	,
(	58075	)	,
(	58111	)	,
(	58148	)	,
(	58184	)	,
(	58221	)	,
(	58257	)	,
(	58294	)	,
(	58330	)	,
(	58367	)	,
(	58403	)	,
(	58439	)	,
(	58476	)	,
(	58512	)	,
(	58549	)	,
(	58585	)	,
(	58622	)	,
(	58658	)	,
(	58695	)	,
(	58731	)	,
(	58768	)	,
(	58804	)	,
(	58840	)	,
(	58877	)	,
(	58913	)	,
(	58950	)	,
(	58986	)	,
(	59023	)	,
(	59059	)	,
(	59096	)	,
(	59132	)	,
(	59168	)	,
(	59205	)	,
(	59241	)	,
(	59278	)	,
(	59314	)	,
(	59351	)	,
(	59387	)	,
(	59424	)	,
(	59460	)	,
(	59497	)	,
(	59533	)	,
(	59569	)	,
(	59606	)	,
(	59642	)	,
(	59679	)	,
(	59715	)	,
(	59752	)	,
(	59788	)	,
(	59825	)	,
(	59861	)	,
(	59898	)	,
(	59934	)	,
(	59970	)	,
(	60007	)	,
(	60043	)	,
(	60080	)	,
(	60116	)	,
(	60153	)	,
(	60189	)	,
(	60226	)	,
(	60262	)	,
(	60298	)	,
(	60335	)	,
(	60371	)	,
(	60408	)	,
(	60444	)	,
(	60481	)	,
(	60517	)	,
(	60554	)	,
(	60590	)	,
(	60627	)	,
(	60663	)	,
(	60699	)	,
(	60736	)	,
(	60772	)	,
(	60809	)	,
(	60845	)	,
(	60882	)	,
(	60918	)	,
(	60955	)	,
(	60991	)	,
(	61028	)	,
(	61064	)	,
(	61100	)	,
(	61137	)	,
(	61173	)	,
(	61210	)	,
(	61246	)	,
(	61283	)	,
(	61319	)	,
(	61356	)	,
(	61392	)	,
(	61429	)	,
(	61465	)	,
(	61501	)	,
(	61538	)	,
(	61574	)	,
(	61611	)	,
(	61647	)	,
(	61684	)	,
(	61720	)	,
(	61757	)	,
(	61793	)	,
(	61829	)	,
(	61866	)	,
(	61902	)	,
(	61939	)	,
(	61975	)	,
(	62012	)	,
(	62048	)	,
(	62085	)	,
(	62121	)	,
(	62158	)	,
(	62194	)	,
(	62230	)	,
(	62267	)	,
(	62303	)	,
(	62340	)	,
(	62376	)	,
(	62413	)	,
(	62449	)	,
(	62486	)	,
(	62522	)	,
(	62559	)	,
(	62595	)	,
(	62631	)	,
(	62668	)	,
(	62704	)	,
(	62741	)	,
(	62777	)	,
(	62814	)	,
(	62850	)	,
(	62887	)	,
(	62923	)	,
(	62959	)	,
(	62996	)	,
(	63032	)	,
(	63069	)	,
(	63105	)	,
(	63142	)	,
(	63178	)	,
(	63215	)	,
(	63251	)	,
(	63288	)	,
(	63324	)	,
(	63360	)	,
(	63397	)	,
(	63433	)	,
(	63470	)	,
(	63506	)	,
(	63543	)	,
(	63579	)	,
(	63616	)	,
(	63652	)	,
(	63689	)	,
(	63725	)	,
(	63761	)	,
(	63798	)	,
(	63834	)	,
(	63871	)	,
(	63907	)	,
(	63944	)	,
(	63980	)	,
(	64017	)	,
(	64053	)	,
(	64090	)	,
(	64126	)	,
(	64162	)	,
(	64199	)	,
(	64235	)	,
(	64272	)	,
(	64308	)	,
(	64345	)	,
(	64381	)	,
(	64418	)	,
(	64454	)	,
(	64490	)	,
(	64527	)	,
(	64563	)	,
(	64600	)	,
(	64636	)	,
(	64673	)	,
(	64709	)	,
(	64746	)	,
(	64782	)	,
(	64819	)	,
(	64855	)	,
(	64891	)	,
(	64928	)	,
(	64964	)	,
(	65001	)	,  -- max distance = max period  = min frequnecy 
(	65037	)	,
(	65074	)	,
(	65110	)	,
(	65147	)	,
(	65183	)	,
(	65220	)	,
(	65256	)	,
(	65292	)	,
(	65329	)	,
(	65365	)	,
(	65402	)	,
(	65438	)	,
(	65475	)	,
(	65511	)	,
(	65548	)	,
(	65584	)	,
(	65620	)	,
(	65657	)	,
(	65693	)	,
(	65730	)	,
(	65766	)	,
(	65803	)	,
(	65839	)	,
(	65876	)	,
(	65912	)	,
(	65949	)	,
(	65985	)	,
(	66021	)	,
(	66058	)	,
(	66094	)	,
(	66131	)	,
(	66167	)	,
(	66204	)	,
(	66240	)	,
(	66277	)	,
(	66313	)	,
(	66350	)	,
(	66386	)	,
(	66422	)	,
(	66459	)	,
(	66495	)	,
(	66532	)	,
(	66568	)	,
(	66605	)	,
(	66641	)	,
(	66678	)	,
(	66714	)	,
(	66750	)	,
(	66787	)	,
(	66823	)	,
(	66860	)	,
(	66896	)	,
(	66933	)	,
(	66969	)	,
(	67006	)	,
(	67042	)	,
(	67079	)	,
(	67115	)	,
(	67151	)	,
(	67188	)	,
(	67224	)	,
(	67261	)	,
(	67297	)	,
(	67334	)	,
(	67370	)	,
(	67407	)	,
(	67443	)	,
(	67480	)	,
(	67516	)	,
(	67552	)	,
(	67589	)	,
(	67625	)	,
(	67662	)	,
(	67698	)	,
(	67735	)	,
(	67771	)	,
(	67808	)	,
(	67844	)	,
(	67881	)	,
(	67917	)	,
(	67953	)	,
(	67990	)	,
(	68026	)	,
(	68063	)	,
(	68099	)	,
(	68136	)	,
(	68172	)	,
(	68209	)	,
(	68245	)	,
(	68281	)	,
(	68318	)	,
(	68354	)	,
(	68391	)	,
(	68427	)	,
(	68464	)	,
(	68500	)	,
(	68537	)	,
(	68573	)	,
(	68610	)	,
(	68646	)	,
(	68682	)	,
(	68719	)	,
(	68755	)	,
(	68792	)	,
(	68828	)	,
(	68865	)	,
(	68901	)	,
(	68938	)	,
(	68974	)	,
(	69011	)	,
(	69047	)	,
(	69083	)	,
(	69120	)	,
(	69156	)	,
(	69193	)	,
(	69229	)	,
(	69266	)	,
(	69302	)	,
(	69339	)	,
(	69375	)	,
(	69411	)	,
(	69448	)	,
(	69484	)	,
(	69521	)	,
(	69557	)	,
(	69594	)	,
(	69630	)	,
(	69667	)	,
(	69703	)	,
(	69740	)	,
(	69776	)	,
(	69812	)	,
(	69849	)	,
(	69885	)	,
(	69922	)	,
(	69958	)	,
(	69995	)	,
(	70031	)	,
(	70068	)	,
(	70104	)	,
(	70141	)	,
(	70177	)	,
(	70213	)	,
(	70250	)	,
(	70286	)	,
(	70323	)	,
(	70359	)	,
(	70396	)	,
(	70432	)	,
(	70469	)	,
(	70505	)	,
(	70542	)	,
(	70578	)	,
(	70614	)	,
(	70651	)	,
(	70687	)	,
(	70724	)	,
(	70760	)	,
(	70797	)	,
(	70833	)	,
(	70870	)	,
(	70906	)	,
(	70942	)	,
(	70979	)	,
(	71015	)	,
(	71052	)	,
(	71088	)	,
(	71125	)	,
(	71161	)	,
(	71198	)	,
(	71234	)	,
(	71271	)	,
(	71307	)	,
(	71343	)	,
(	71380	)	,
(	71416	)	,
(	71453	)	,
(	71489	)	,
(	71526	)	,
(	71562	)	,
(	71599	)	,
(	71635	)	,
(	71672	)	,
(	71708	)	,
(	71744	)	,
(	71781	)	,
(	71817	)	,
(	71854	)	,
(	71890	)	,
(	71927	)	,
(	71963	)	,
(	72000	)	,
(	72036	)	,
(	72072	)	,
(	72109	)	,
(	72145	)	,
(	72182	)	,
(	72218	)	,
(	72255	)	,
(	72291	)	,
(	72328	)	,
(	72364	)	,
(	72401	)	,
(	72437	)	,
(	72473	)	,
(	72510	)	,
(	72546	)	,
(	72583	)	,
(	72619	)	,
(	72656	)	,
(	72692	)	,
(	72729	)	,
(	72765	)	,
(	72802	)	,
(	72838	)	,
(	72874	)	,
(	72911	)	,
(	72947	)	,
(	72984	)	,
(	73020	)	,
(	73057	)	,
(	73093	)	,
(	73130	)	,
(	73166	)	,
(	73203	)	,
(	73239	)	,
(	73275	)	,
(	73312	)	,
(	73348	)	,
(	73385	)	,
(	73421	)	,
(	73458	)	,
(	73494	)	,
(	73531	)	,
(	73567	)	,
(	73603	)	,
(	73640	)	,
(	73676	)	,
(	73713	)	,
(	73749	)	,
(	73786	)	,
(	73822	)	,
(	73859	)	,
(	73895	)	,
(	73932	)	,
(	73968	)	,
(	74004	)	,
(	74041	)	,
(	74077	)	,
(	74114	)	,
(	74150	)	,
(	74187	)	,
(	74223	)	,
(	74260	)	,
(	74296	)	,
(	74333	)	,
(	74369	)	,
(	74405	)	,
(	74442	)	,
(	74478	)	,
(	74515	)	,
(	74551	)	,
(	74588	)	,
(	74624	)	,
(	74661	)	,
(	74697	)	,
(	74733	)	,
(	74770	)	,
(	74806	)	,
(	74843	)	,
(	74879	)	,
(	74916	)	,
(	74952	)	,
(	74989	)	,
(	75025	)	,
(	75062	)	,
(	75098	)	,
(	75134	)	,
(	75171	)	,
(	75207	)	,
(	75244	)	,
(	75280	)	,
(	75317	)	,
(	75353	)	,
(	75390	)	,
(	75426	)	,
(	75463	)	,
(	75499	)	,
(	75535	)	,
(	75572	)	,
(	75608	)	,
(	75645	)	,
(	75681	)	,
(	75718	)	,
(	75754	)	,
(	75791	)	,
(	75827	)	,
(	75863	)	,
(	75900	)	,
(	75936	)	,
(	75973	)	,
(	76009	)	,
(	76046	)	,
(	76082	)	,
(	76119	)	,
(	76155	)	,
(	76192	)	,
(	76228	)	,
(	76264	)	,
(	76301	)	,
(	76337	)	,
(	76374	)	,
(	76410	)	,
(	76447	)	,
(	76483	)	,
(	76520	)	,
(	76556	)	,
(	76593	)	,
(	76629	)	,
(	76665	)	,
(	76702	)	,
(	76738	)	,
(	76775	)	,
(	76811	)	,
(	76848	)	,
(	76884	)	,
(	76921	)	,
(	76957	)	,
(	76994	)	,
(	77030	)	,
(	77066	)	,
(	77103	)	,
(	77139	)	,
(	77176	)	,
(	77212	)	,
(	77249	)	,
(	77285	)	,
(	77322	)	,
(	77358	)	,
(	77394	)	,
(	77431	)	,
(	77467	)	,
(	77504	)	,
(	77540	)	,
(	77577	)	,
(	77613	)	,
(	77650	)	,
(	77686	)	,
(	77723	)	,
(	77759	)	,
(	77795	)	,
(	77832	)	,
(	77868	)	,
(	77905	)	,
(	77941	)	,
(	77978	)	,
(	78014	)	,
(	78051	)	,
(	78087	)	,
(	78124	)	,
(	78160	)	,
(	78196	)	,
(	78233	)	,
(	78269	)	,
(	78306	)	,
(	78342	)	,
(	78379	)	,
(	78415	)	,
(	78452	)	,
(	78488	)	,
(	78524	)	,
(	78561	)	,
(	78597	)	,
(	78634	)	,
(	78670	)	,
(	78707	)	,
(	78743	)	,
(	78780	)	,
(	78816	)	,
(	78853	)	,
(	78889	)	,
(	78925	)	,
(	78962	)	,
(	78998	)	,
(	79035	)	,
(	79071	)	,
(	79108	)	,
(	79144	)	,
(	79181	)	,
(	79217	)	,
(	79254	)	,
(	79290	)	,
(	79326	)	,
(	79363	)	,
(	79399	)	,
(	79436	)	,
(	79472	)	,
(	79509	)	,
(	79545	)	,
(	79582	)	,
(	79618	)	,
(	79655	)	,
(	79691	)	,
(	79727	)	,
(	79764	)	,
(	79800	)	,
(	79837	)	,
(	79873	)	,
(	79910	)	,
(	79946	)	,
(	79983	)	,
(	80019	)	,
(	80055	)	,
(	80092	)	,
(	80128	)	,
(	80165	)	,
(	80201	)	,
(	80238	)	,
(	80274	)	,
(	80311	)	,
(	80347	)	,
(	80384	)	,
(	80420	)	,
(	80456	)	,
(	80493	)	,
(	80529	)	,
(	80566	)	,
(	80602	)	,
(	80639	)	,
(	80675	)	,
(	80712	)	,
(	80748	)	,
(	80785	)	,
(	80821	)	,
(	80857	)	,
(	80894	)	,
(	80930	)	,
(	80967	)	,
(	81003	)	,
(	81040	)	,
(	81076	)	,
(	81113	)	,
(	81149	)	,
(	81185	)	,
(	81222	)	,
(	81258	)	,
(	81295	)	,
(	81331	)	,
(	81368	)	,
(	81404	)	,
(	81441	)	,
(	81477	)	,
(	81514	)	,
(	81550	)	,
(	81586	)	,
(	81623	)	,
(	81659	)	,
(	81696	)	,
(	81732	)	,
(	81769	)	,
(	81805	)	,
(	81842	)	,
(	81878	)	,
(	81915	)	,
(	81951	)	,
(	81987	)	,
(	82024	)	,
(	82060	)	,
(	82097	)	,
(	82133	)	,
(	82170	)	,
(	82206	)	,
(	82243	)	,
(	82279	)	,
(	82316	)	,
(	82352	)	,
(	82388	)	,
(	82425	)	,
(	82461	)	,
(	82498	)	,
(	82534	)	,
(	82571	)	,
(	82607	)	,
(	82644	)	,
(	82680	)	,
(	82716	)	,
(	82753	)	,
(	82789	)	,
(	82826	)	,
(	82862	)	,
(	82899	)	,
(	82935	)	,
(	82972	)	,
(	83008	)	,
(	83045	)	,
(	83081	)	,
(	83117	)	,
(	83154	)	,
(	83190	)	,
(	83227	)	,
(	83263	)	,
(	83300	)	,
(	83336	)	,
(	83373	)	,
(	83409	)	,
(	83446	)	,
(	83482	)	,
(	83518	)	,
(	83555	)	,
(	83591	)	,
(	83628	)	,
(	83664	)	,
(	83701	)	,
(	83737	)	,
(	83774	)	,
(	83810	)	,
(	83846	)	,
(	83883	)	,
(	83919	)	,
(	83956	)	,
(	83992	)	,
(	84029	)	,
(	84065	)	,
(	84102	)	,
(	84138	)	,
(	84175	)	,
(	84211	)	,
(	84247	)	,
(	84284	)	,
(	84320	)	,
(	84357	)	,
(	84393	)	,
(	84430	)	,
(	84466	)	,
(	84503	)	,
(	84539	)	,
(	84576	)	,
(	84612	)	,
(	84648	)	,
(	84685	)	,
(	84721	)	,
(	84758	)	,
(	84794	)	,
(	84831	)	,
(	84867	)	,
(	84904	)	,
(	84940	)	,
(	84976	)	,
(	85013	)	,
(	85049	)	,
(	85086	)	,
(	85122	)	,
(	85159	)	,
(	85195	)	,
(	85232	)	,
(	85268	)	,
(	85305	)	,
(	85341	)	,
(	85377	)	,
(	85414	)	,
(	85450	)	,
(	85487	)	,
(	85523	)	,
(	85560	)	,
(	85596	)	,
(	85633	)	,
(	85669	)	,
(	85706	)	,
(	85742	)	,
(	85778	)	,
(	85815	)	,
(	85851	)	,
(	85888	)	,
(	85924	)	,
(	85961	)	,
(	85997	)	,
(	86034	)	,
(	86070	)	,
(	86107	)	,
(	86143	)	,
(	86179	)	,
(	86216	)	,
(	86252	)	,
(	86289	)	,
(	86325	)	,
(	86362	)	,
(	86398	)	,
(	86435	)	,
(	86471	)	,
(	86507	)	,
(	86544	)	,
(	86580	)	,
(	86617	)	,
(	86653	)	,
(	86690	)	,
(	86726	)	,
(	86763	)	,
(	86799	)	,
(	86836	)	,
(	86872	)	,
(	86908	)	,
(	86945	)	,
(	86981	)	,
(	87018	)	,
(	87054	)	,
(	87091	)	,
(	87127	)	,
(	87164	)	,
(	87200	)	,
(	87237	)	,
(	87273	)	,
(	87309	)	,
(	87346	)	,
(	87382	)	,
(	87419	)	,
(	87455	)	,
(	87492	)	,
(	87528	)	,
(	87565	)	,
(	87601	)	,
(	87637	)	,
(	87674	)	,
(	87710	)	,
(	87747	)	,
(	87783	)	,
(	87820	)	,
(	87856	)	,
(	87893	)	,
(	87929	)	,
(	87966	)	,
(	88002	)	,
(	88038	)	,
(	88075	)	,
(	88111	)	,
(	88148	)	,
(	88184	)	,
(	88221	)	,
(	88257	)	,
(	88294	)	,
(	88330	)	,
(	88367	)	,
(	88403	)	,
(	88439	)	,
(	88476	)	,
(	88512	)	,
(	88549	)	,
(	88585	)	,
(	88622	)	,
(	88658	)	,
(	88695	)	,
(	88731	)	,
(	88768	)	,
(	88804	)	,
(	88840	)	,
(	88877	)	,
(	88913	)	,
(	88950	)	,
(	88986	)	,
(	89023	)	,
(	89059	)	,
(	89096	)	,
(	89132	)	,
(	89168	)	,
(	89205	)	,
(	89241	)	,
(	89278	)	,
(	89314	)	,
(	89351	)	,
(	89387	)	,
(	89424	)	,
(	89460	)	,
(	89497	)	,
(	89533	)	,
(	89569	)	,
(	89606	)	,
(	89642	)	,
(	89679	)	,
(	89715	)	,
(	89752	)	,
(	89788	)	,
(	89825	)	,
(	89861	)	,
(	89898	)	,
(	89934	)	,
(	89970	)	,
(	90007	)	,
(	90043	)	,
(	90080	)	,
(	90116	)	,
(	90153	)	,
(	90189	)	,
(	90226	)	,
(	90262	)	,
(	90298	)	,
(	90335	)	,
(	90371	)	,
(	90408	)	,
(	90444	)	,
(	90481	)	,
(	90517	)	,
(	90554	)	,
(	90590	)	,
(	90627	)	,
(	90663	)	,
(	90699	)	,
(	90736	)	,
(	90772	)	,
(	90809	)	,
(	90845	)	,
(	90882	)	,
(	90918	)	,
(	90955	)	,
(	90991	)	,
(	91028	)	,
(	91064	)	,
(	91100	)	,
(	91137	)	,
(	91173	)	,
(	91210	)	,
(	91246	)	,
(	91283	)	,
(	91319	)	,
(	91356	)	,
(	91392	)	,
(	91429	)	,
(	91465	)	,
(	91501	)	,
(	91538	)	,
(	91574	)	,
(	91611	)	,
(	91647	)	,
(	91684	)	,
(	91720	)	,
(	91757	)	,
(	91793	)	,
(	91829	)	,
(	91866	)	,
(	91902	)	,
(	91939	)	,
(	91975	)	,
(	92012	)	,
(	92048	)	,
(	92085	)	,
(	92121	)	,
(	92158	)	,
(	92194	)	,
(	92230	)	,
(	92267	)	,
(	92303	)	,
(	92340	)	,
(	92376	)	,
(	92413	)	,
(	92449	)	,
(	92486	)	,
(	92522	)	,
(	92559	)	,
(	92595	)	,
(	92631	)	,
(	92668	)	,
(	92704	)	,
(	92741	)	,
(	92777	)	,
(	92814	)	,
(	92850	)	,
(	92887	)	,
(	92923	)	,
(	92959	)	,
(	92996	)	,
(	93032	)	,
(	93069	)	,
(	93105	)	,
(	93142	)	,
(	93178	)	,
(	93215	)	,
(	93251	)	,
(	93288	)	,
(	93324	)	,
(	93360	)	,
(	93397	)	,
(	93433	)	,
(	93470	)	,
(	93506	)	,
(	93543	)	,
(	93579	)	,
(	93616	)	,
(	93652	)	,
(	93689	)	,
(	93725	)	,
(	93761	)	,
(	93798	)	,
(	93834	)	,
(	93871	)	,
(	93907	)	,
(	93944	)	,
(	93980	)	,
(	94017	)	,
(	94053	)	,
(	94089	)	,
(	94126	)	,
(	94162	)	,
(	94199	)	,
(	94235	)	,
(	94272	)	,
(	94308	)	,
(	94345	)	,
(	94381	)	,
(	94418	)	,
(	94454	)	,
(	94490	)	,
(	94527	)	,
(	94563	)	,
(	94600	)	,
(	94636	)	,
(	94673	)	,
(	94709	)	,
(	94746	)	,
(	94782	)	,
(	94819	)	,
(	94855	)	,
(	94891	)	,
(	94928	)	,
(	94964	)	,
(	95001	)	,
(	95037	)	,
(	95074	)	,
(	95110	)	,
(	95147	)	,
(	95183	)	,
(	95220	)	,
(	95256	)	,
(	95292	)	,
(	95329	)	,
(	95365	)	,
(	95402	)	,
(	95438	)	,
(	95475	)	,
(	95511	)	,
(	95548	)	,
(	95584	)	,
(	95620	)	,
(	95657	)	,
(	95693	)	,
(	95730	)	,
(	95766	)	,
(	95803	)	,
(	95839	)	,
(	95876	)	,
(	95912	)	,
(	95949	)	,
(	95985	)	,
(	96021	)	,
(	96058	)	,
(	96094	)	,
(	96131	)	,
(	96167	)	,
(	96204	)	,
(	96240	)	,
(	96277	)	,
(	96313	)	,
(	96350	)	,
(	96386	)	,
(	96422	)	,
(	96459	)	,
(	96495	)	,
(	96532	)	,
(	96568	)	,
(	96605	)	,
(	96641	)	,
(	96678	)	,
(	96714	)	,
(	96750	)	,
(	96787	)	,
(	96823	)	,
(	96860	)	,
(	96896	)	,
(	96933	)	,
(	96969	)	,
(	97006	)	,
(	97042	)	,
(	97079	)	,
(	97115	)	,
(	97151	)	,
(	97188	)	,
(	97224	)	,
(	97261	)	,
(	97297	)	,
(	97334	)	,
(	97370	)	,
(	97407	)	,
(	97443	)	,
(	97480	)	,
(	97516	)	,
(	97552	)	,
(	97589	)	,
(	97625	)	,
(	97662	)	,
(	97698	)	,
(	97735	)	,
(	97771	)	,
(	97808	)	,
(	97844	)	,
(	97881	)	,
(	97917	)	,
(	97953	)	,
(	97990	)	,
(	98026	)	,
(	98063	)	,
(	98099	)	,
(	98136	)	,
(	98172	)	,
(	98209	)	,
(	98245	)	,
(	98281	)	,
(	98318	)	,
(	98354	)	,
(	98391	)	,
(	98427	)	,
(	98464	)	,
(	98500	)	,
(	98537	)	,
(	98573	)	,
(	98610	)	,
(	98646	)	,
(	98682	)	,
(	98719	)	,
(	98755	)	,
(	98792	)	,
(	98828	)	,
(	98865	)	,
(	98901	)	,
(	98938	)	,
(	98974	)	,
(	99011	)	,
(	99047	)	,
(	99083	)	,
(	99120	)	,
(	99156	)	,
(	99193	)	,
(	99229	)	,
(	99266	)	,
(	99302	)	,
(	99339	)	,
(	99375	)	,
(	99411	)	,
(	99448	)	,
(	99484	)	,
(	99521	)	,
(	99557	)	,
(	99594	)	,
(	99630	)	,
(	99667	)	,
(	99703	)	,
(	99740	)	,
(	99776	)	,
(	99812	)	,
(	99849	)	,
(	99885	)	,
(	99922	)	,
(	99958	)	,
(	99995	)	,
(	100031	)	,
(	100068	)	,
(	100104	)	,
(	100141	)	,
(	100177	)	,
(	100213	)	,
(	100250	)	,
(	100286	)	,
(	100323	)	,
(	100359	)	,
(	100396	)	,
(	100432	)	,
(	100469	)	,
(	100505	)	,
(	100542	)	,
(	100578	)	,
(	100614	)	,
(	100651	)	,
(	100687	)	,
(	100724	)	,
(	100760	)	,
(	100797	)	,
(	100833	)	,
(	100870	)	,
(	100906	)	,
(	100942	)	,
(	100979	)	,
(	101015	)	,
(	101052	)	,
(	101088	)	,
(	101125	)	,
(	101161	)	,
(	101198	)	,
(	101234	)	,
(	101271	)	,
(	101307	)	,
(	101343	)	,
(	101380	)	,
(	101416	)	,
(	101453	)	,
(	101489	)	,
(	101526	)	,
(	101562	)	,
(	101599	)	,
(	101635	)	,
(	101672	)	,
(	101708	)	,
(	101744	)	,
(	101781	)	,
(	101817	)	,
(	101854	)	,
(	101890	)	,
(	101927	)	,
(	101963	)	,
(	102000	)	,
(	102036	)	,
(	102072	)	,
(	102109	)	,
(	102145	)	,
(	102182	)	,
(	102218	)	,
(	102255	)	,
(	102291	)	,
(	102328	)	,
(	102364	)	,
(	102401	)	,
(	102437	)	,
(	102473	)	,
(	102510	)	,
(	102546	)	,
(	102583	)	,
(	102619	)	,
(	102656	)	,
(	102692	)	,
(	102729	)	,
(	102765	)	,
(	102802	)	,
(	102838	)	,
(	102874	)	,
(	102911	)	,
(	102947	)	,
(	102984	)	,
(	103020	)	,
(	103057	)	,
(	103093	)	,
(	103130	)	,
(	103166	)	,
(	103202	)	,
(	103239	)	,
(	103275	)	,
(	103312	)	,
(	103348	)	,
(	103385	)	,
(	103421	)	,
(	103458	)	,
(	103494	)	,
(	103531	)	,
(	103567	)	,
(	103603	)	,
(	103640	)	,
(	103676	)	,
(	103713	)	,
(	103749	)	,
(	103786	)	,
(	103822	)	,
(	103859	)	,
(	103895	)	,
(	103932	)	,
(	103968	)	,
(	104004	)	,
(	104041	)	,
(	104077	)	,
(	104114	)	,
(	104150	)	,
(	104187	)	,
(	104223	)	,
(	104260	)	,
(	104296	)	,
(	104333	)	,
(	104369	)	,
(	104405	)	,
(	104442	)	,
(	104478	)	,
(	104515	)	,
(	104551	)	,
(	104588	)	,
(	104624	)	,
(	104661	)	,
(	104697	)	,
(	104733	)	,
(	104770	)	,
(	104806	)	,
(	104843	)	,
(	104879	)	,
(	104916	)	,
(	104952	)	,
(	104989	)	,
(	105025	)	,
(	105062	)	,
(	105098	)	,
(	105134	)	,
(	105171	)	,
(	105207	)	,
(	105244	)	,
(	105280	)	,
(	105317	)	,
(	105353	)	,
(	105390	)	,
(	105426	)	,
(	105463	)	,
(	105499	)	,
(	105535	)	,
(	105572	)	,
(	105608	)	,
(	105645	)	,
(	105681	)	,
(	105718	)	,
(	105754	)	,
(	105791	)	,
(	105827	)	,
(	105863	)	,
(	105900	)	,
(	105936	)	,
(	105973	)	,
(	106009	)	,
(	106046	)	,
(	106082	)	,
(	106119	)	,
(	106155	)	,
(	106192	)	,
(	106228	)	,
(	106264	)	,
(	106301	)	,
(	106337	)	,
(	106374	)	,
(	106410	)	,
(	106447	)	,
(	106483	)	,
(	106520	)	,
(	106556	)	,
(	106593	)	,
(	106629	)	,
(	106665	)	,
(	106702	)	,
(	106738	)	,
(	106775	)	,
(	106811	)	,
(	106848	)	,
(	106884	)	,
(	106921	)	,
(	106957	)	,
(	106994	)	,
(	107030	)	,
(	107066	)	,
(	107103	)	,
(	107139	)	,
(	107176	)	,
(	107212	)	,
(	107249	)	,
(	107285	)	,
(	107322	)	,
(	107358	)	,
(	107394	)	,
(	107431	)	,
(	107467	)	,
(	107504	)	,
(	107540	)	,
(	107577	)	,
(	107613	)	,
(	107650	)	,
(	107686	)	,
(	107723	)	,
(	107759	)	,
(	107795	)	,
(	107832	)	,
(	107868	)	,
(	107905	)	,
(	107941	)	,
(	107978	)	,
(	108014	)	,
(	108051	)	,
(	108087	)	,
(	108124	)	,
(	108160	)	,
(	108196	)	,
(	108233	)	,
(	108269	)	,
(	108306	)	,
(	108342	)	,
(	108379	)	,
(	108415	)	,
(	108452	)	,
(	108488	)	,
(	108524	)	,
(	108561	)	,
(	108597	)	,
(	108634	)	,
(	108670	)	,
(	108707	)	,
(	108743	)	,
(	108780	)	,
(	108816	)	,
(	108853	)	,
(	108889	)	,
(	108925	)	,
(	108962	)	,
(	108998	)	,
(	109035	)	,
(	109071	)	,
(	109108	)	,
(	109144	)	,
(	109181	)	,
(	109217	)	,
(	109254	)	,
(	109290	)	,
(	109326	)	,
(	109363	)	,
(	109399	)	,
(	109436	)	,
(	109472	)	,
(	109509	)	,
(	109545	)	,
(	109582	)	,
(	109618	)	,
(	109655	)	,
(	109691	)	,
(	109727	)	,
(	109764	)	,
(	109800	)	,
(	109837	)	,
(	109873	)	,
(	109910	)	,
(	109946	)	,
(	109983	)	,
(	110019	)	,
(	110055	)	,
(	110092	)	,
(	110128	)	,
(	110165	)	,
(	110201	)	,
(	110238	)	,
(	110274	)	,
(	110311	)	,
(	110347	)	,
(	110384	)	,
(	110420	)	,
(	110456	)	,
(	110493	)	,
(	110529	)	,
(	110566	)	,
(	110602	)	,
(	110639	)	,
(	110675	)	,
(	110712	)	,
(	110748	)	,
(	110785	)	,
(	110821	)	,
(	110857	)	,
(	110894	)	,
(	110930	)	,
(	110967	)	,
(	111003	)	,
(	111040	)	,
(	111076	)	,
(	111113	)	,
(	111149	)	,
(	111185	)	,
(	111222	)	,
(	111258	)	,
(	111295	)	,
(	111331	)	,
(	111368	)	,
(	111404	)	,
(	111441	)	,
(	111477	)	,
(	111514	)	,
(	111550	)	,
(	111586	)	,
(	111623	)	,
(	111659	)	,
(	111696	)	,
(	111732	)	,
(	111769	)	,
(	111805	)	,
(	111842	)	,
(	111878	)	,
(	111915	)	,
(	111951	)	,
(	111987	)	,
(	112024	)	,
(	112060	)	,
(	112097	)	,
(	112133	)	,
(	112170	)	,
(	112206	)	,
(	112243	)	,
(	112279	)	,
(	112315	)	,
(	112352	)	,
(	112388	)	,
(	112425	)	,
(	112461	)	,
(	112498	)	,
(	112534	)	,
(	112571	)	,
(	112607	)	,
(	112644	)	,
(	112680	)	,
(	112716	)	,
(	112753	)	,
(	112789	)	,
(	112826	)	,
(	112862	)	,
(	112899	)	,
(	112935	)	,
(	112972	)	,
(	113008	)	,
(	113045	)	,
(	113081	)	,
(	113117	)	,
(	113154	)	,
(	113190	)	,
(	113227	)	,
(	113263	)	,
(	113300	)	,
(	113336	)	,
(	113373	)	,
(	113409	)	,
(	113446	)	,
(	113482	)	,
(	113518	)	,
(	113555	)	,
(	113591	)	,
(	113628	)	,
(	113664	)	,
(	113701	)	,
(	113737	)	,
(	113774	)	,
(	113810	)	,
(	113846	)	,
(	113883	)	,
(	113919	)	,
(	113956	)	,
(	113992	)	,
(	114029	)	,
(	114065	)	,
(	114102	)	,
(	114138	)	,
(	114175	)	,
(	114211	)	,
(	114247	)	,
(	114284	)	,
(	114320	)	,
(	114357	)	,
(	114393	)	,
(	114430	)	,
(	114466	)	,
(	114503	)	,
(	114539	)	,
(	114576	)	,
(	114612	)	,
(	114648	)	,
(	114685	)	,
(	114721	)	,
(	114758	)	,
(	114794	)	,
(	114831	)	,
(	114867	)	,
(	114904	)	,
(	114940	)	,
(	114976	)	,
(	115013	)	,
(	115049	)	,
(	115086	)	,
(	115122	)	,
(	115159	)	,
(	115195	)	,
(	115232	)	,
(	115268	)	,
(	115305	)	,
(	115341	)	,
(	115377	)	,
(	115414	)	,
(	115450	)	,
(	115487	)	,
(	115523	)	,
(	115560	)	,
(	115596	)	,
(	115633	)	,
(	115669	)	,
(	115706	)	,
(	115742	)	,
(	115778	)	,
(	115815	)	,
(	115851	)	,
(	115888	)	,
(	115924	)	,
(	115961	)	,
(	115997	)	,
(	116034	)	,
(	116070	)	,
(	116107	)	,
(	116143	)	,
(	116179	)	,
(	116216	)	,
(	116252	)	,
(	116289	)	,
(	116325	)	,
(	116362	)	,
(	116398	)	,
(	116435	)	,
(	116471	)	,
(	116507	)	,
(	116544	)	,
(	116580	)	,
(	116617	)	,
(	116653	)	,
(	116690	)	,
(	116726	)	,
(	116763	)	,
(	116799	)	,
(	116836	)	,
(	116872	)	,
(	116908	)	,
(	116945	)	,
(	116981	)	,
(	117018	)	,
(	117054	)	,
(	117091	)	,
(	117127	)	,
(	117164	)	,
(	117200	)	,
(	117237	)	,
(	117273	)	,
(	117309	)	,
(	117346	)	,
(	117382	)	,
(	117419	)	,
(	117455	)	,
(	117492	)	,
(	117528	)	,
(	117565	)	,
(	117601	)	,
(	117637	)	,
(	117674	)	,
(	117710	)	,
(	117747	)	,
(	117783	)	,
(	117820	)	,
(	117856	)	,
(	117893	)	,
(	117929	)	,
(	117966	)	,
(	118002	)	,
(	118038	)	,
(	118075	)	,
(	118111	)	,
(	118148	)	,
(	118184	)	,
(	118221	)	,
(	118257	)	,
(	118294	)	,
(	118330	)	,
(	118367	)	,
(	118403	)	,
(	118439	)	,
(	118476	)	,
(	118512	)	,
(	118549	)	,
(	118585	)	,
(	118622	)	,
(	118658	)	,
(	118695	)	,
(	118731	)	,
(	118768	)	,
(	118804	)	,
(	118840	)	,
(	118877	)	,
(	118913	)	,
(	118950	)	,
(	118986	)	,
(	119023	)	,
(	119059	)	,
(	119096	)	,
(	119132	)	,
(	119168	)	,
(	119205	)	,
(	119241	)	,
(	119278	)	,
(	119314	)	,
(	119351	)	,
(	119387	)	,
(	119424	)	,
(	119460	)	,
(	119497	)	,
(	119533	)	,
(	119569	)	,
(	119606	)	,
(	119642	)	,
(	119679	)	,
(	119715	)	,
(	119752	)	,
(	119788	)	,
(	119825	)	,
(	119861	)	,
(	119898	)	,
(	119934	)	,
(	119970	)	,
(	120007	)	,
(	120043	)	,
(	120080	)	,
(	120116	)	,
(	120153	)	,
(	120189	)	,
(	120226	)	,
(	120262	)	,
(	120298	)	,
(	120335	)	,
(	120371	)	,
(	120408	)	,
(	120444	)	,
(	120481	)	,
(	120517	)	,
(	120554	)	,
(	120590	)	,
(	120627	)	,
(	120663	)	,
(	120699	)	,
(	120736	)	,
(	120772	)	,
(	120809	)	,
(	120845	)	,
(	120882	)	,
(	120918	)	,
(	120955	)	,
(	120991	)	,
(	121028	)	,
(	121064	)	,
(	121100	)	,
(	121137	)	,
(	121173	)	,
(	121210	)	,
(	121246	)	,
(	121283	)	,
(	121319	)	,
(	121356	)	,
(	121392	)	,
(	121428	)	,
(	121465	)	,
(	121501	)	,
(	121538	)	,
(	121574	)	,
(	121611	)	,
(	121647	)	,
(	121684	)	,
(	121720	)	,
(	121757	)	,
(	121793	)	,
(	121829	)	,
(	121866	)	,
(	121902	)	,
(	121939	)	,
(	121975	)	,
(	122012	)	,
(	122048	)	,
(	122085	)	,
(	122121	)	,
(	122158	)	,
(	122194	)	,
(	122230	)	,
(	122267	)	,
(	122303	)	,
(	122340	)	,
(	122376	)	,
(	122413	)	,
(	122449	)	,
(	122486	)	,
(	122522	)	,
(	122559	)	,
(	122595	)	,
(	122631	)	,
(	122668	)	,
(	122704	)	,
(	122741	)	,
(	122777	)	,
(	122814	)	,
(	122850	)	,
(	122887	)	,
(	122923	)	,
(	122959	)	,
(	122996	)	,
(	123032	)	,
(	123069	)	,
(	123105	)	,
(	123142	)	,
(	123178	)	,
(	123215	)	,
(	123251	)	,
(	123288	)	,
(	123324	)	,
(	123360	)	,
(	123397	)	,
(	123433	)	,
(	123470	)	,
(	123506	)	,
(	123543	)	,
(	123579	)	,
(	123616	)	,
(	123652	)	,
(	123689	)	,
(	123725	)	,
(	123761	)	,
(	123798	)	,
(	123834	)	,
(	123871	)	,
(	123907	)	,
(	123944	)	,
(	123980	)	,
(	124017	)	,
(	124053	)	,
(	124089	)	,
(	124126	)	,
(	124162	)	,
(	124199	)	,
(	124235	)	,
(	124272	)	,
(	124308	)	,
(	124345	)	,
(	124381	)	,
(	124418	)	,
(	124454	)	,
(	124490	)	,
(	124527	)	,
(	124563	)	,
(	124600	)	,
(	124636	)	,
(	124673	)	,
(	124709	)	,
(	124746	)	,
(	124782	)	,
(	124819	)	,
(	124855	)	,
(	124891	)	,
(	124928	)	,
(	124964	)	,
(	125001	)	,
(	125037	)	,
(	125074	)	,
(	125110	)	,
(	125147	)	,
(	125183	)	,
(	125220	)	,
(	125256	)	,
(	125292	)	,
(	125329	)	,
(	125365	)	,
(	125402	)	,
(	125438	)	,
(	125475	)	,
(	125511	)	,
(	125548	)	,
(	125584	)	,
(	125620	)	,
(	125657	)	,
(	125693	)	,
(	125730	)	,
(	125766	)	,
(	125803	)	,
(	125839	)	,
(	125876	)	,
(	125912	)	,
(	125949	)	,
(	125985	)	,
(	126021	)	,
(	126058	)	,
(	126094	)	,
(	126131	)	,
(	126167	)	,
(	126204	)	,
(	126240	)	,
(	126277	)	,
(	126313	)	,
(	126350	)	,
(	126386	)	,
(	126422	)	,
(	126459	)	,
(	126495	)	,
(	126532	)	,
(	126568	)	,
(	126605	)	,
(	126641	)	,
(	126678	)	,
(	126714	)	,
(	126750	)	,
(	126787	)	,
(	126823	)	,
(	126860	)	,
(	126896	)	,
(	126933	)	,
(	126969	)	,
(	127006	)	,
(	127042	)	,
(	127079	)	,
(	127115	)	,
(	127151	)	,
(	127188	)	,
(	127224	)	,
(	127261	)	,
(	127297	)	,
(	127334	)	,
(	127370	)	,
(	127407	)	,
(	127443	)	,
(	127480	)	,
(	127516	)	,
(	127552	)	,
(	127589	)	,
(	127625	)	,
(	127662	)	,
(	127698	)	,
(	127735	)	,
(	127771	)	,
(	127808	)	,
(	127844	)	,
(	127881	)	,
(	127917	)	,
(	127953	)	,
(	127990	)	,
(	128026	)	,
(	128063	)	,
(	128099	)	,
(	128136	)	,
(	128172	)	,
(	128209	)	,
(	128245	)	,
(	128281	)	,
(	128318	)	,
(	128354	)	,
(	128391	)	,
(	128427	)	,
(	128464	)	,
(	128500	)	,
(	128537	)	,
(	128573	)	,
(	128610	)	,
(	128646	)	,
(	128682	)	,
(	128719	)	,
(	128755	)	,
(	128792	)	,
(	128828	)	,
(	128865	)	,
(	128901	)	,
(	128938	)	,
(	128974	)	,
(	129011	)	,
(	129047	)	,
(	129083	)	,
(	129120	)	,
(	129156	)	,
(	129193	)	,
(	129229	)	,
(	129266	)	,
(	129302	)	,
(	129339	)	,
(	129375	)	,
(	129411	)	,
(	129448	)	,
(	129484	)	,
(	129521	)	,
(	129557	)	,
(	129594	)	,
(	129630	)	,
(	129667	)	,
(	129703	)	,
(	129740	)	,
(	129776	)	,
(	129812	)	,
(	129849	)	,
(	129885	)	,
(	129922	)	,
(	129958	)	,
(	129995	)	,
(	130031	)	,
(	130068	)	,
(	130104	)	,
(	130141	)	,
(	130177	)	,
(	130213	)	,
(	130250	)	,
(	130286	)	,
(	130323	)	,
(	130359	)	,
(	130396	)	,
(	130432	)	,
(	130469	)	,
(	130505	)	,
(	130541	)	,
(	130578	)	,
(	130614	)	,
(	130651	)	,
(	130687	)	,
(	130724	)	,
(	130760	)	,
(	130797	)	,
(	130833	)	,
(	130870	)	,
(	130906	)	,
(	130942	)	,
(	130979	)	,
(	131015	)	,
(	131052	)	,
(	131088	)	,
(	131125	)	,
(	131161	)	,
(	131198	)	,
(	131234	)	,
(	131271	)	,
(	131307	)	,
(	131343	)	,
(	131380	)	,
(	131416	)	,
(	131453	)	,
(	131489	)	,
(	131526	)	,
(	131562	)	,
(	131599	)	,
(	131635	)	,
(	131672	)	,
(	131708	)	,
(	131744	)	,
(	131781	)	,
(	131817	)	,
(	131854	)	,
(	131890	)	,
(	131927	)	,
(	131963	)	,
(	132000	)	,
(	132036	)	,
(	132072	)	,
(	132109	)	,
(	132145	)	,
(	132182	)	,
(	132218	)	,
(	132255	)	,
(	132291	)	,
(	132328	)	,
(	132364	)	,
(	132401	)	,
(	132437	)	,
(	132473	)	,
(	132510	)	,
(	132546	)	,
(	132583	)	,
(	132619	)	,
(	132656	)	,
(	132692	)	,
(	132729	)	,
(	132765	)	,
(	132802	)	,
(	132838	)	,
(	132874	)	,
(	132911	)	,
(	132947	)	,
(	132984	)	,
(	133020	)	,
(	133057	)	,
(	133093	)	,
(	133130	)	,
(	133166	)	,
(	133202	)	,
(	133239	)	,
(	133275	)	,
(	133312	)	,
(	133348	)	,
(	133385	)	,
(	133421	)	,
(	133458	)	,
(	133494	)	,
(	133531	)	,
(	133567	)	,
(	133603	)	,
(	133640	)	,
(	133676	)	,
(	133713	)	,
(	133749	)	,
(	133786	)	,
(	133822	)	,
(	133859	)	,
(	133895	)	,
(	133932	)	,
(	133968	)	,
(	134004	)	,
(	134041	)	,
(	134077	)	,
(	134114	)	,
(	134150	)	,
(	134187	)	,
(	134223	)	,
(	134260	)	,
(	134296	)	,
(	134333	)	,
(	134369	)	,
(	134405	)	,
(	134442	)	,
(	134478	)	,
(	134515	)	,
(	134551	)	,
(	134588	)	,
(	134624	)	,
(	134661	)	,
(	134697	)	,
(	134733	)	,
(	134770	)	,
(	134806	)	,
(	134843	)	,
(	134879	)	,
(	134916	)	,
(	134952	)	,
(	134989	)	,
(	135025	)	,
(	135062	)	,
(	135098	)	,
(	135134	)	,
(	135171	)	,
(	135207	)	,
(	135244	)	,
(	135280	)	,
(	135317	)	,
(	135353	)	,
(	135390	)	,
(	135426	)	,
(	135463	)	,
(	135499	)	,
(	135535	)	,
(	135572	)	,
(	135608	)	,
(	135645	)	,
(	135681	)	,
(	135718	)	,
(	135754	)	,
(	135791	)	,
(	135827	)	,
(	135863	)	,
(	135900	)	,
(	135936	)	,
(	135973	)	,
(	136009	)	,
(	136046	)	,
(	136082	)	,
(	136119	)	,
(	136155	)	,
(	136192	)	,
(	136228	)	,
(	136264	)	,
(	136301	)	,
(	136337	)	,
(	136374	)	,
(	136410	)	,
(	136447	)	,
(	136483	)	,
(	136520	)	,
(	136556	)	,
(	136593	)	,
(	136629	)	,
(	136665	)	,
(	136702	)	,
(	136738	)	,
(	136775	)	,
(	136811	)	,
(	136848	)	,
(	136884	)	,
(	136921	)	,
(	136957	)	,
(	136994	)	,
(	137030	)	,
(	137066	)	,
(	137103	)	,
(	137139	)	,
(	137176	)	,
(	137212	)	,
(	137249	)	,
(	137285	)	,
(	137322	)	,
(	137358	)	,
(	137394	)	,
(	137431	)	,
(	137467	)	,
(	137504	)	,
(	137540	)	,
(	137577	)	,
(	137613	)	,
(	137650	)	,
(	137686	)	,
(	137723	)	,
(	137759	)	,
(	137795	)	,
(	137832	)	,
(	137868	)	,
(	137905	)	,
(	137941	)	,
(	137978	)	,
(	138014	)	,
(	138051	)	,
(	138087	)	,
(	138124	)	,
(	138160	)	,
(	138196	)	,
(	138233	)	,
(	138269	)	,
(	138306	)	,
(	138342	)	,
(	138379	)	,
(	138415	)	,
(	138452	)	,
(	138488	)	,
(	138524	)	,
(	138561	)	,
(	138597	)	,
(	138634	)	,
(	138670	)	,
(	138707	)	,
(	138743	)	,
(	138780	)	,
(	138816	)	,
(	138853	)	,
(	138889	)	,
(	138925	)	,
(	138962	)	,
(	138998	)	,
(	139035	)	,
(	139071	)	,
(	139108	)	,
(	139144	)	,
(	139181	)	,
(	139217	)	,
(	139254	)	,
(	139290	)	,
(	139326	)	,
(	139363	)	,
(	139399	)	,
(	139436	)	,
(	139472	)	,
(	139509	)	,
(	139545	)	,
(	139582	)	,
(	139618	)	,
(	139654	)	,
(	139691	)	,
(	139727	)	,
(	139764	)	,
(	139800	)	,
(	139837	)	,
(	139873	)	,
(	139910	)	,
(	139946	)	,
(	139983	)	,
(	140019	)	,
(	140055	)	,
(	140092	)	,
(	140128	)	,
(	140165	)	,
(	140201	)	,
(	140238	)	,
(	140274	)	,
(	140311	)	,
(	140347	)	,
(	140384	)	,
(	140420	)	,
(	140456	)	,
(	140493	)	,
(	140529	)	,
(	140566	)	,
(	140602	)	,
(	140639	)	,
(	140675	)	,
(	140712	)	,
(	140748	)	,
(	140785	)	,
(	140821	)	,
(	140857	)	,
(	140894	)	,
(	140930	)	,
(	140967	)	,
(	141003	)	,
(	141040	)	,
(	141076	)	,
(	141113	)	,
(	141149	)	,
(	141185	)	,
(	141222	)	,
(	141258	)	,
(	141295	)	,
(	141331	)	,
(	141368	)	, 
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	,
(	141368	)	

);

end package LUT_flashing_pkg;